module TLMonitor(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_a_bits_corrupt,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [2:0]  io_in_c_bits_size,
  input  [6:0]  io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [6:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input         io_in_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_86 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_2 = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_3 = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_4 = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_5 = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_lo = mask_acc_2 | mask_size_2 & mask_eq_6; // @[Misc.scala 214:29]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_hi = mask_acc_2 | mask_size_2 & mask_eq_7; // @[Misc.scala 214:29]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_lo = mask_acc_3 | mask_size_2 & mask_eq_8; // @[Misc.scala 214:29]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_hi = mask_acc_3 | mask_size_2 & mask_eq_9; // @[Misc.scala 214:29]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_lo = mask_acc_4 | mask_size_2 & mask_eq_10; // @[Misc.scala 214:29]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_hi = mask_acc_4 | mask_size_2 & mask_eq_11; // @[Misc.scala 214:29]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_lo = mask_acc_5 | mask_size_2 & mask_eq_12; // @[Misc.scala 214:29]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_hi = mask_acc_5 | mask_size_2 & mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire [31:0] _T_180 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_181 = {1'b0,$signed(_T_180)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_183 = $signed(_T_181) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_184 = $signed(_T_183) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_185 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_186 = {1'b0,$signed(_T_185)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_188 = $signed(_T_186) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_189 = $signed(_T_188) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_190 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_191 = {1'b0,$signed(_T_190)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_193 = $signed(_T_191) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_194 = $signed(_T_193) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_195 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_196 = {1'b0,$signed(_T_195)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_198 = $signed(_T_196) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_199 = $signed(_T_198) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_200 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_201 = {1'b0,$signed(_T_200)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_203 = $signed(_T_201) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_204 = $signed(_T_203) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_211 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_214 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_215 = {1'b0,$signed(_T_214)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_217 = $signed(_T_215) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_218 = $signed(_T_217) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_219 = _T_211 & _T_218; // @[Parameters.scala 670:56]
  wire  _T_222 = source_ok & _T_219; // @[Monitor.scala 82:72]
  wire  _T_277 = _source_ok_T_1 & _T_211; // @[Mux.scala 27:72]
  wire  _T_330 = _T_218 | _T_184 | _T_189 | _T_194 | _T_199 | _T_204; // @[Parameters.scala 671:42]
  wire  _T_333 = _T_277 & _T_330; // @[Monitor.scala 83:78]
  wire  _T_347 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [7:0] _T_351 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_352 = _T_351 == 8'h0; // @[Monitor.scala 88:31]
  wire  _T_356 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18]
  wire  _T_360 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_593 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_606 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_709 = _T_211 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_720 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_724 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_732 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_834 = source_ok & _T_709; // @[Monitor.scala 115:71]
  wire  _T_852 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [7:0] _T_968 = ~mask; // @[Monitor.scala 127:33]
  wire [7:0] _T_969 = io_in_a_bits_mask & _T_968; // @[Monitor.scala 127:31]
  wire  _T_970 = _T_969 == 8'h0; // @[Monitor.scala 127:40]
  wire  _T_974 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_1088 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_1096 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_1210 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_1218 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1332 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1344 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1348 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1352 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27]
  wire  _T_1356 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_1360 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1364 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1368 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1379 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_1383 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_1396 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1416 = _T_1364 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1425 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1442 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1460 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _source_ok_T_109 = io_in_c_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_115 = io_in_c_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_121 = io_in_c_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_127 = io_in_c_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_133 = io_in_c_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_139 = io_in_c_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_145 = io_in_c_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_151 = io_in_c_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_2 = _source_ok_T_109 | _source_ok_T_115 | _source_ok_T_121 | _source_ok_T_127 | _source_ok_T_133 |
    _source_ok_T_139 | _source_ok_T_145 | _source_ok_T_151; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_7 = 13'h3f << io_in_c_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask_2 = ~_is_aligned_mask_T_7[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_87 = {{26'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T_2 = io_in_c_bits_address & _GEN_87; // @[Edges.scala 20:16]
  wire  is_aligned_2 = _is_aligned_T_2 == 32'h0; // @[Edges.scala 20:24]
  wire [31:0] _address_ok_T_34 = io_in_c_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_35 = {1'b0,$signed(_address_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_37 = $signed(_address_ok_T_35) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_38 = $signed(_address_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_39 = io_in_c_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_40 = {1'b0,$signed(_address_ok_T_39)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_42 = $signed(_address_ok_T_40) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_43 = $signed(_address_ok_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_44 = io_in_c_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_45 = {1'b0,$signed(_address_ok_T_44)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_47 = $signed(_address_ok_T_45) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_48 = $signed(_address_ok_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_49 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_50 = {1'b0,$signed(_address_ok_T_49)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_52 = $signed(_address_ok_T_50) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_53 = $signed(_address_ok_T_52) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_54 = io_in_c_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_55 = {1'b0,$signed(_address_ok_T_54)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_57 = $signed(_address_ok_T_55) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_58 = $signed(_address_ok_T_57) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _address_ok_T_62 = _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 | _address_ok_T_58; // @[Parameters.scala 598:92]
  wire [31:0] _address_ok_T_63 = io_in_c_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_64 = {1'b0,$signed(_address_ok_T_63)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_66 = $signed(_address_ok_T_64) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_67 = $signed(_address_ok_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  wire  address_ok_1 = _address_ok_T_62 | _address_ok_T_67; // @[Parameters.scala 622:64]
  wire  _T_2230 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  wire  _T_2237 = io_in_c_bits_size >= 3'h3; // @[Monitor.scala 245:30]
  wire  _T_2244 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  wire  _T_2252 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  wire  _T_2270 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  wire  _T_2363 = io_in_c_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_2371 = _T_2363 & _address_ok_T_67; // @[Parameters.scala 670:56]
  wire  _T_2374 = source_ok_2 & _T_2371; // @[Monitor.scala 260:78]
  wire  _T_2429 = _source_ok_T_109 & _T_2363; // @[Mux.scala 27:72]
  wire  _T_2482 = _address_ok_T_67 | _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 |
    _address_ok_T_58; // @[Parameters.scala 671:42]
  wire  _T_2485 = _T_2429 & _T_2482; // @[Monitor.scala 261:78]
  wire  _T_2507 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  wire  _T_2740 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  wire  _T_2750 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  wire  _T_2758 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  wire  _T_2772 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  wire  sink_ok_1 = io_in_e_bits_sink < 1'h1; // @[Monitor.scala 364:31]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [6:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_2794 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_2795 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_2799 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_2803 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_2807 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_2811 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [6:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_2818 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_2819 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_2823 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_2827 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_2831 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_2839 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  wire  _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  wire [2:0] c_first_beats1_decode = is_aligned_mask_2[5:3]; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  reg [2:0] c_first_counter; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1 = c_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  c_first = c_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [2:0] size_3; // @[Monitor.scala 514:22]
  reg [6:0] source_3; // @[Monitor.scala 515:22]
  reg [31:0] address_2; // @[Monitor.scala 516:22]
  wire  _T_2870 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  wire  _T_2871 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  wire  _T_2875 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  wire  _T_2879 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  wire  _T_2883 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  wire  _T_2887 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  reg [127:0] inflight; // @[Monitor.scala 611:27]
  reg [511:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [511:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  wire [8:0] _GEN_88 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [9:0] _a_opcode_lookup_T = {{1'd0}, _GEN_88}; // @[Monitor.scala 634:69]
  wire [511:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [511:0] _GEN_89 = {{496'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_89; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[511:1]}; // @[Monitor.scala 634:152]
  wire [511:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [511:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 638:91]
  wire [511:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[511:1]}; // @[Monitor.scala 638:144]
  wire  _T_2893 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [127:0] _a_set_wo_ready_T = 128'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_2896 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [8:0] _GEN_94 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [9:0] _a_opcodes_set_T = {{1'd0}, _GEN_94}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [1026:0] _GEN_95 = {{1023'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [1026:0] _a_opcodes_set_T_1 = _GEN_95 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [1026:0] _GEN_97 = {{1023'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [1026:0] _a_sizes_set_T_1 = _GEN_97 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [127:0] _T_2898 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_2900 = ~_T_2898[0]; // @[Monitor.scala 658:17]
  wire [127:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [1026:0] _GEN_31 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [1026:0] _GEN_32 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_2904 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_2906 = ~_T_1348; // @[Monitor.scala 671:74]
  wire  _T_2907 = io_in_d_valid & d_first_1 & ~_T_1348; // @[Monitor.scala 671:71]
  wire [127:0] _d_clr_wo_ready_T = 128'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1348 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [1038:0] _GEN_99 = {{1023'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [1038:0] _d_opcodes_clr_T_5 = _GEN_99 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [127:0] d_clr = _d_first_T & d_first_1 & _T_2906 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [1038:0] _GEN_35 = _d_first_T & d_first_1 & _T_2906 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_2893 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [127:0] _T_2917 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_2919 = _T_2917[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_2924 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_2925 = io_in_d_bits_opcode == _GEN_44 | _T_2924; // @[Monitor.scala 685:77]
  wire  _T_2929 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_2936 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_2937 = io_in_d_bits_opcode == _GEN_60 | _T_2936; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_102 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_2941 = _GEN_102 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_2951 = _T_2904 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_2906; // @[Monitor.scala 694:116]
  wire  _T_2952 = ~io_in_d_ready; // @[Monitor.scala 695:15]
  wire  _T_2953 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_2960 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [127:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [127:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [127:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [511:0] a_opcodes_set = _GEN_31[511:0];
  wire [511:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [511:0] d_opcodes_clr = _GEN_35[511:0];
  wire [511:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [511:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [511:0] a_sizes_set = _GEN_32[511:0];
  wire [511:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [511:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_2969 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [127:0] inflight_1; // @[Monitor.scala 723:35]
  reg [511:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [2:0] c_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1_1 = c_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  c_first_1 = c_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25]
  wire [511:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [511:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 747:93]
  wire [511:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[511:1]}; // @[Monitor.scala 747:146]
  wire  _T_2979 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  _T_2980 = io_in_c_valid & c_first_1 & _T_2979; // @[Monitor.scala 756:37]
  wire [127:0] _c_set_wo_ready_T = 128'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] c_set_wo_ready = io_in_c_valid & c_first_1 & _T_2979 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 756:71 Monitor.scala 757:22]
  wire  _T_2986 = _c_first_T & c_first_1 & _T_2979; // @[Monitor.scala 760:38]
  wire [3:0] _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  wire [3:0] _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 4'h1; // @[Monitor.scala 763:59]
  wire [8:0] _GEN_109 = {io_in_c_bits_source, 2'h0}; // @[Monitor.scala 764:79]
  wire [9:0] _c_opcodes_set_T = {{1'd0}, _GEN_109}; // @[Monitor.scala 764:79]
  wire [3:0] c_sizes_set_interm = _c_first_T & c_first_1 & _T_2979 ? _c_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 760:72 Monitor.scala 763:28]
  wire [1026:0] _GEN_112 = {{1023'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  wire [1026:0] _c_sizes_set_T_1 = _GEN_112 << _c_opcodes_set_T; // @[Monitor.scala 765:52]
  wire [127:0] _T_2987 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  wire  _T_2989 = ~_T_2987[0]; // @[Monitor.scala 766:17]
  wire [127:0] c_set = _c_first_T & c_first_1 & _T_2979 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 760:72 Monitor.scala 761:28]
  wire [1026:0] _GEN_77 = _c_first_T & c_first_1 & _T_2979 ? _c_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 760:72 Monitor.scala 765:28]
  wire  _T_2993 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  wire  _T_2995 = io_in_d_valid & d_first_2 & _T_1348; // @[Monitor.scala 779:71]
  wire [127:0] d_clr_wo_ready_1 = io_in_d_valid & d_first_2 & _T_1348 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 779:89 Monitor.scala 780:22]
  wire [127:0] d_clr_1 = _d_first_T & d_first_2 & _T_1348 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [1038:0] _GEN_80 = _d_first_T & d_first_2 & _T_1348 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire  _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1 = _T_2980 & io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:88]
  wire [127:0] _T_3003 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire  _T_3005 = _T_3003[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  wire  _T_3009 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_3013 = _GEN_102 == c_size_lookup; // @[Monitor.scala 795:36]
  wire  _T_3022 = _T_2993 & c_first_1 & io_in_c_valid & _same_cycle_resp_T_8 & _T_1348; // @[Monitor.scala 799:116]
  wire  _T_3024 = _T_2952 | io_in_c_ready; // @[Monitor.scala 800:32]
  wire  _T_3028 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  wire  _T_3029 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  wire [127:0] _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  wire [127:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [127:0] _inflight_T_5 = _inflight_T_3 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [511:0] d_opcodes_clr_1 = _GEN_80[511:0];
  wire [511:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [511:0] c_sizes_set = _GEN_77[511:0];
  wire [511:0] _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  wire [511:0] _inflight_sizes_T_5 = _inflight_sizes_T_3 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_3038 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [2:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_3 = d_first_counter_3 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 3'h0; // @[Edges.scala 230:25]
  wire  _T_3050 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_3051 = _d_first_T & d_first_3 & _T_3050; // @[Monitor.scala 829:38]
  wire  _T_3054 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = _d_first_T & d_first_3 & _T_3050 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  _T_3058 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _e_clr_T = 2'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  wire  d_set = _GEN_84[0];
  wire  _T_3062 = (d_set | inflight_2) >> io_in_e_bits_sink; // @[Monitor.scala 837:35]
  wire [1:0] _GEN_85 = _T_3058 ? _e_clr_T : 2'h0; // @[Monitor.scala 835:73 Monitor.scala 836:13]
  wire  e_clr = _GEN_85[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 3'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      opcode_3 <= io_in_c_bits_opcode; // @[Monitor.scala 525:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      param_3 <= io_in_c_bits_param; // @[Monitor.scala 526:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      size_3 <= io_in_c_bits_size; // @[Monitor.scala 527:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      source_3 <= io_in_c_bits_source; // @[Monitor.scala 528:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      address_2 <= io_in_c_bits_address; // @[Monitor.scala 529:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 128'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 512'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 512'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 128'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 512'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first_1) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 3'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_c_first_T | _d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= (inflight_2 | d_set) & ~e_clr; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 3'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_356 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_356 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_356 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1088 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1088 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(_T_1210 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(_T_1210 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1096 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(_T_1332 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(_T_1332 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(_T_356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1218 & ~(_T_356 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1344 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1344 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(_T_1360 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(_T_1360 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(_T_1364 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1348 & ~(_T_1364 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(_T_1379 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(_T_1379 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(_T_1383 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(_T_1383 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(_T_1360 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1368 & ~(_T_1360 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(_T_1379 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(_T_1379 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(_T_1383 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(_T_1383 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(_T_1416 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1396 & ~(_T_1416 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1425 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1425 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1425 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1425 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1425 & ~(_T_1360 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1425 & ~(_T_1360 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1442 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1442 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1442 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1442 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1442 & ~(_T_1416 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1442 & ~(_T_1416 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1460 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1460 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1460 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1460 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1460 & ~(_T_1360 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1460 & ~(_T_1360 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(_T_2237 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(_T_2237 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(_T_2244 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2230 & ~(_T_2244 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(_T_2237 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(_T_2237 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(_T_2244 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2252 & ~(_T_2244 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(_T_2374 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(_T_2374 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(_T_2485 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(_T_2485 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(_T_2237 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(_T_2237 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(_T_2244 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid report param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2270 & ~(_T_2244 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(_T_2374 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(_T_2374 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(_T_2485 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(_T_2485 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(_T_2237 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(_T_2237 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(_T_2244 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2507 & ~(_T_2244 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2740 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2740 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2740 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2740 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2740 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2740 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2740 & ~(_T_2750 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2740 & ~(_T_2750 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2758 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2758 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2758 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2758 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2758 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2758 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2758 & ~(_T_2750 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2758 & ~(_T_2750 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2772 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2772 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2772 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2772 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2772 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2772 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2772 & ~(_T_2750 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2772 & ~(_T_2750 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channels carries invalid sink ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2794 & ~(_T_2795 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2794 & ~(_T_2795 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2794 & ~(_T_2799 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2794 & ~(_T_2799 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2794 & ~(_T_2803 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2794 & ~(_T_2803 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2794 & ~(_T_2807 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2794 & ~(_T_2807 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2794 & ~(_T_2811 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2794 & ~(_T_2811 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2818 & ~(_T_2819 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2818 & ~(_T_2819 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2818 & ~(_T_2823 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2818 & ~(_T_2823 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2818 & ~(_T_2827 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2818 & ~(_T_2827 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2818 & ~(_T_2831 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2818 & ~(_T_2831 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2818 & ~(_T_2839 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2818 & ~(_T_2839 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2870 & ~(_T_2871 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2870 & ~(_T_2871 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2870 & ~(_T_2875 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2870 & ~(_T_2875 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2870 & ~(_T_2879 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2870 & ~(_T_2879 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2870 & ~(_T_2883 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2870 & ~(_T_2883 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2870 & ~(_T_2887 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2870 & ~(_T_2887 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2896 & ~(_T_2900 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2896 & ~(_T_2900 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2907 & ~(_T_2919 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2907 & ~(_T_2919 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2907 & same_cycle_resp & ~(_T_2925 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2907 & same_cycle_resp & ~(_T_2925 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2907 & same_cycle_resp & ~(_T_2929 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2907 & same_cycle_resp & ~(_T_2929 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2907 & ~same_cycle_resp & ~(_T_2937 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2907 & ~same_cycle_resp & ~(_T_2937 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2907 & ~same_cycle_resp & ~(_T_2941 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2907 & ~same_cycle_resp & ~(_T_2941 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2951 & ~(_T_2953 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2951 & ~(_T_2953 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2960 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2960 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2969 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2969 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2986 & ~(_T_2989 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel re-used a source ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2986 & ~(_T_2989 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2995 & ~(_T_3005 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2995 & ~(_T_3005 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2995 & same_cycle_resp_1 & ~(_T_3009 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2995 & same_cycle_resp_1 & ~(_T_3009 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2995 & ~same_cycle_resp_1 & ~(_T_3013 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2995 & ~same_cycle_resp_1 & ~(_T_3013 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3022 & ~(_T_3024 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3022 & ~(_T_3024 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3028 & ~(_T_3029 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3028 & ~(_T_3029 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_3038 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_3038 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3051 & ~(_T_3054 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3051 & ~(_T_3054 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3058 & ~(_T_3062 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:8)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3058 & ~(_T_3062 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  c_first_counter = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  opcode_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  param_3 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  size_3 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  source_3 = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  address_2 = _RAND_17[31:0];
  _RAND_18 = {4{`RANDOM}};
  inflight = _RAND_18[127:0];
  _RAND_19 = {16{`RANDOM}};
  inflight_opcodes = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  inflight_sizes = _RAND_20[511:0];
  _RAND_21 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  watchdog = _RAND_23[31:0];
  _RAND_24 = {4{`RANDOM}};
  inflight_1 = _RAND_24[127:0];
  _RAND_25 = {16{`RANDOM}};
  inflight_sizes_1 = _RAND_25[511:0];
  _RAND_26 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  watchdog_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inflight_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_30[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_a_bits_corrupt,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [2:0]  auto_in_c_bits_size,
  input  [6:0]  auto_in_c_bits_source,
  input  [31:0] auto_in_c_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  output        auto_in_e_ready,
  input         auto_in_e_valid,
  input         auto_in_e_bits_sink,
  input         auto_out_1_a_ready,
  output        auto_out_1_a_valid,
  output [2:0]  auto_out_1_a_bits_opcode,
  output [2:0]  auto_out_1_a_bits_param,
  output [2:0]  auto_out_1_a_bits_size,
  output [6:0]  auto_out_1_a_bits_source,
  output [12:0] auto_out_1_a_bits_address,
  output [7:0]  auto_out_1_a_bits_mask,
  output        auto_out_1_a_bits_corrupt,
  input         auto_out_1_c_ready,
  output        auto_out_1_c_valid,
  output [2:0]  auto_out_1_c_bits_opcode,
  output [2:0]  auto_out_1_c_bits_param,
  output [2:0]  auto_out_1_c_bits_size,
  output [6:0]  auto_out_1_c_bits_source,
  output [12:0] auto_out_1_c_bits_address,
  output        auto_out_1_d_ready,
  input         auto_out_1_d_valid,
  input  [2:0]  auto_out_1_d_bits_opcode,
  input  [1:0]  auto_out_1_d_bits_param,
  input  [2:0]  auto_out_1_d_bits_size,
  input  [6:0]  auto_out_1_d_bits_source,
  input         auto_out_1_d_bits_denied,
  input         auto_out_1_d_bits_corrupt,
  output        auto_out_1_e_valid,
  input         auto_out_0_a_ready,
  output        auto_out_0_a_valid,
  output [2:0]  auto_out_0_a_bits_opcode,
  output [2:0]  auto_out_0_a_bits_param,
  output [2:0]  auto_out_0_a_bits_size,
  output [6:0]  auto_out_0_a_bits_source,
  output [31:0] auto_out_0_a_bits_address,
  output [7:0]  auto_out_0_a_bits_mask,
  output [63:0] auto_out_0_a_bits_data,
  output        auto_out_0_a_bits_corrupt,
  output        auto_out_0_d_ready,
  input         auto_out_0_d_valid,
  input  [2:0]  auto_out_0_d_bits_opcode,
  input  [2:0]  auto_out_0_d_bits_size,
  input  [6:0]  auto_out_0_d_bits_source,
  input         auto_out_0_d_bits_denied,
  input  [63:0] auto_out_0_d_bits_data,
  input         auto_out_0_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_bits_sink; // @[Nodes.scala 24:25]
  reg [2:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 3'h0; // @[Arbiter.scala 88:28]
  wire [1:0] readys_filter_lo = {auto_out_1_d_valid,auto_out_0_d_valid}; // @[Cat.scala 30:58]
  reg [1:0] readys_mask; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 24:30]
  wire [1:0] readys_filter_hi = readys_filter_lo & _readys_filter_T; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter = {readys_filter_hi,auto_out_1_d_valid,auto_out_0_d_valid}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_1 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_1; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_2 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready = _GEN_2 | _readys_unready_T_4; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  wire  readys_0 = readys_readys[0]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_0 = readys_0 & auto_out_0_d_valid; // @[Arbiter.scala 97:79]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire [6:0] _T_36 = muxStateEarly_0 ? auto_out_0_d_bits_source : 7'h0; // @[Mux.scala 27:72]
  wire  readys_1 = readys_readys[1]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_1 = readys_1 & auto_out_1_d_valid; // @[Arbiter.scala 97:79]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire [6:0] _T_37 = muxStateEarly_1 ? auto_out_1_d_bits_source : 7'h0; // @[Mux.scala 27:72]
  wire [31:0] _requestAIO_T = auto_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_1 = {1'b0,$signed(_requestAIO_T)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_3 = $signed(_requestAIO_T_1) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_4 = $signed(_requestAIO_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_5 = auto_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_6 = {1'b0,$signed(_requestAIO_T_5)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_8 = $signed(_requestAIO_T_6) & 33'she0000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_9 = $signed(_requestAIO_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_10 = auto_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_11 = {1'b0,$signed(_requestAIO_T_10)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_13 = $signed(_requestAIO_T_11) & 33'shc0000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_14 = $signed(_requestAIO_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_15 = auto_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_16 = {1'b0,$signed(_requestAIO_T_15)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_18 = $signed(_requestAIO_T_16) & 33'shc0000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_19 = $signed(_requestAIO_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_20 = auto_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_21 = {1'b0,$signed(_requestAIO_T_20)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_23 = $signed(_requestAIO_T_21) & 33'she0000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_24 = $signed(_requestAIO_T_23) == 33'sh0; // @[Parameters.scala 137:67]
  wire  requestAIO_0_0 = _requestAIO_T_4 | _requestAIO_T_9 | _requestAIO_T_14 | _requestAIO_T_19 | _requestAIO_T_24; // @[Xbar.scala 363:92]
  wire [32:0] _requestAIO_T_30 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_32 = $signed(_requestAIO_T_30) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_1 = $signed(_requestAIO_T_32) == 33'sh0; // @[Parameters.scala 137:67]
  wire  requestEIO_0_1 = ~auto_in_e_bits_sink; // @[Parameters.scala 46:9]
  wire [12:0] _beatsDO_decode_T_1 = 13'h3f << auto_out_0_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_3 = ~_beatsDO_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode = _beatsDO_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata = auto_out_0_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] beatsDO_0 = beatsDO_opdata ? beatsDO_decode : 3'h0; // @[Edges.scala 220:14]
  wire [12:0] _beatsDO_decode_T_5 = 13'h3f << auto_out_1_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_7 = ~_beatsDO_decode_T_5[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode_1 = _beatsDO_decode_T_7[5:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata_1 = auto_out_1_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] beatsDO_1 = beatsDO_opdata_1 ? beatsDO_decode_1 : 3'h0; // @[Edges.scala 220:14]
  wire  latch = idle & auto_in_d_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _readys_mask_T = readys_readys & readys_filter_lo; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 244:43]
  wire  _prefixOR_T = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 104:53]
  wire  _T_10 = auto_out_0_d_valid | auto_out_1_d_valid; // @[Arbiter.scala 107:36]
  wire  _T_11 = ~(auto_out_0_d_valid | auto_out_1_d_valid); // @[Arbiter.scala 107:15]
  wire [2:0] maskedBeats_0 = earlyWinner_0 ? beatsDO_0 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_1 = earlyWinner_1 ? beatsDO_1 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] initBeats = maskedBeats_0 | maskedBeats_1; // @[Arbiter.scala 112:44]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & auto_out_0_d_valid | state_1 & auto_out_1_d_valid; // @[Mux.scala 27:72]
  wire  sink_ACancel_5_earlyValid = idle ? _T_10 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_5_earlyValid; // @[ReadyValidCancel.scala 50:33]
  wire [2:0] _GEN_3 = {{2'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [2:0] _beatsLeft_T_4 = beatsLeft - _GEN_3; // @[Arbiter.scala 113:52]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire [2:0] _T_39 = muxStateEarly_0 ? auto_out_0_d_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_40 = muxStateEarly_1 ? auto_out_1_d_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_45 = muxStateEarly_0 ? auto_out_0_d_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_46 = muxStateEarly_1 ? auto_out_1_d_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  TLMonitor monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_c_ready(monitor_io_in_c_ready),
    .io_in_c_valid(monitor_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_io_in_c_bits_address),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),
    .io_in_e_ready(monitor_io_in_e_ready),
    .io_in_e_valid(monitor_io_in_e_valid),
    .io_in_e_bits_sink(monitor_io_in_e_bits_sink)
  );
  assign auto_in_a_ready = requestAIO_0_0 & auto_out_0_a_ready | requestAIO_0_1 & auto_out_1_a_ready; // @[Mux.scala 27:72]
  assign auto_in_c_ready = auto_out_1_c_ready; // @[Mux.scala 27:72]
  assign auto_in_d_valid = idle ? _T_10 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_in_d_bits_opcode = _T_45 | _T_46; // @[Mux.scala 27:72]
  assign auto_in_d_bits_param = muxStateEarly_1 ? auto_out_1_d_bits_param : 2'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_size = _T_39 | _T_40; // @[Mux.scala 27:72]
  assign auto_in_d_bits_source = _T_36 | _T_37; // @[Mux.scala 27:72]
  assign auto_in_d_bits_denied = muxStateEarly_0 & auto_out_0_d_bits_denied | muxStateEarly_1 & auto_out_1_d_bits_denied
    ; // @[Mux.scala 27:72]
  assign auto_in_d_bits_data = muxStateEarly_0 ? auto_out_0_d_bits_data : 64'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_corrupt = muxStateEarly_0 & auto_out_0_d_bits_corrupt | muxStateEarly_1 &
    auto_out_1_d_bits_corrupt; // @[Mux.scala 27:72]
  assign auto_in_e_ready = ~auto_in_e_bits_sink; // @[Parameters.scala 46:9]
  assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1; // @[Xbar.scala 428:50]
  assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_1_a_bits_address = auto_in_a_bits_address[12:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_1_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_c_valid = auto_in_c_valid; // @[ReadyValidCancel.scala 21:38]
  assign auto_out_1_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_c_bits_source = auto_in_c_bits_source; // @[Xbar.scala 259:55]
  assign auto_out_1_c_bits_address = auto_in_c_bits_address[12:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_1_d_ready = auto_in_d_ready & allowed_1; // @[Arbiter.scala 123:31]
  assign auto_out_1_e_valid = auto_in_e_valid & requestEIO_0_1; // @[Xbar.scala 179:40]
  assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0; // @[Xbar.scala 428:50]
  assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_0_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_d_ready = auto_in_d_ready & allowed_0; // @[Arbiter.scala 123:31]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = requestAIO_0_0 & auto_out_0_a_ready | requestAIO_0_1 & auto_out_1_a_ready; // @[Mux.scala 27:72]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_ready = auto_out_1_c_ready; // @[Mux.scala 27:72]
  assign monitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = idle ? _T_10 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign monitor_io_in_d_bits_opcode = _T_45 | _T_46; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_param = muxStateEarly_1 ? auto_out_1_d_bits_param : 2'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_size = _T_39 | _T_40; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_source = _T_36 | _T_37; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_denied = muxStateEarly_0 & auto_out_0_d_bits_denied | muxStateEarly_1 &
    auto_out_1_d_bits_denied; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_corrupt = muxStateEarly_0 & auto_out_0_d_bits_corrupt | muxStateEarly_1 &
    auto_out_1_d_bits_corrupt; // @[Mux.scala 27:72]
  assign monitor_io_in_e_ready = ~auto_in_e_bits_sink; // @[Parameters.scala 46:9]
  assign monitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 3'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin // @[Arbiter.scala 113:23]
      beatsLeft <= initBeats;
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch & |readys_filter_lo) begin // @[Arbiter.scala 27:32]
      readys_mask <= _readys_mask_T_3; // @[Arbiter.scala 28:12]
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin // @[Arbiter.scala 117:30]
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin // @[Arbiter.scala 117:30]
      state_1 <= earlyWinner_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(auto_out_0_d_valid | auto_out_1_d_valid) | _prefixOR_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(auto_out_0_d_valid | auto_out_1_d_valid) | _prefixOR_T | reset)) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_11 | _T_10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_11 | _T_10 | reset)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  readys_mask = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  state_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_1(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [3:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [3:0]  io_in_a_bits_mask,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [3:0]  io_in_d_bits_source,
  input  [5:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = ~io_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | io_in_a_bits_source[3]; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_34 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_60 = 3'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48]
  wire [31:0] _T_62 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_63 = {1'b0,$signed(_T_62)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_65 = $signed(_T_63) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_66 = $signed(_T_65) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_77 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_78 = {1'b0,$signed(_T_77)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_80 = $signed(_T_78) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_81 = $signed(_T_80) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_82 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_83 = {1'b0,$signed(_T_82)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_85 = $signed(_T_83) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_86 = $signed(_T_85) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_90 = _T_66 | _T_71 | _T_76 | _T_81 | _T_86; // @[Parameters.scala 671:42]
  wire  _T_91 = _T_60 & _T_90; // @[Parameters.scala 670:56]
  wire  _T_93 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_96 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_97 = {1'b0,$signed(_T_96)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_99 = $signed(_T_97) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_100 = $signed(_T_99) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_101 = _T_93 & _T_100; // @[Parameters.scala 670:56]
  wire  _T_104 = _T_91 | _T_101; // @[Parameters.scala 672:30]
  wire  _T_105 = source_ok & _T_104; // @[Monitor.scala 82:72]
  wire [32:0] _T_136 = $signed(_T_78) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _T_137 = $signed(_T_136) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_141 = _T_100 | _T_66 | _T_71 | _T_76 | _T_137; // @[Parameters.scala 671:42]
  wire [3:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_163 = _T_162 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_312 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_367 = _T_93 & _T_141; // @[Parameters.scala 670:56]
  wire  _T_382 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_390 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_444 = source_ok & _T_367; // @[Monitor.scala 115:71]
  wire  _T_462 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_530 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_531 = io_in_a_bits_mask & _T_530; // @[Monitor.scala 127:31]
  wire  _T_532 = _T_531 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_536 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_556 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_581 = _T_66 | _T_71 | _T_76 | _T_137; // @[Parameters.scala 671:42]
  wire  _T_582 = _T_556 & _T_581; // @[Parameters.scala 670:56]
  wire  _T_594 = _T_582 | _T_101; // @[Parameters.scala 672:30]
  wire  _T_595 = source_ok & _T_594; // @[Monitor.scala 131:74]
  wire  _T_613 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_690 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_766 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_13 = ~io_in_d_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_13 | io_in_d_bits_source[3]; // @[Parameters.scala 1125:46]
  wire  sink_ok = io_in_d_bits_sink < 6'h21; // @[Monitor.scala 306:31]
  wire  _T_770 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_774 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_778 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_782 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_786 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_790 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_801 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_805 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_818 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_838 = _T_786 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_847 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_864 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_882 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [3:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_912 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_913 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_921 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_925 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_929 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [3:0] source_1; // @[Monitor.scala 538:22]
  reg [5:0] sink; // @[Monitor.scala 539:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_936 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_937 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_941 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_945 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_949 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_953 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29]
  wire  _T_957 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [15:0] inflight; // @[Monitor.scala 611:27]
  reg [63:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [63:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69]
  wire [63:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [63:0] _GEN_73 = {{48'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[63:1]}; // @[Monitor.scala 634:152]
  wire [63:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [63:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91]
  wire [63:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[63:1]}; // @[Monitor.scala 638:144]
  wire  _T_963 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire  _T_966 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [15:0] _T_968 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_970 = ~_T_968[0]; // @[Monitor.scala 658:17]
  wire [15:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [130:0] _GEN_19 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [130:0] _GEN_20 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_974 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_976 = ~_T_770; // @[Monitor.scala 671:74]
  wire  _T_977 = io_in_d_valid & d_first_1 & ~_T_770; // @[Monitor.scala 671:71]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [15:0] d_clr = _d_first_T & d_first_1 & _T_976 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [142:0] _GEN_23 = _d_first_T & d_first_1 & _T_976 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_963 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [15:0] _T_987 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_989 = _T_987[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_994 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39]
  wire  _T_995 = io_in_d_bits_opcode == _GEN_32 | _T_994; // @[Monitor.scala 685:77]
  wire  _T_999 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_1006 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_1007 = io_in_d_bits_opcode == _GEN_48 | _T_1006; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_1011 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_1021 = _T_974 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_976; // @[Monitor.scala 694:116]
  wire  _T_1023 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire [15:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [15:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [15:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [63:0] a_opcodes_set = _GEN_19[63:0];
  wire [63:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [63:0] d_opcodes_clr = _GEN_23[63:0];
  wire [63:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [63:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [63:0] a_sizes_set = _GEN_20[63:0];
  wire [63:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [63:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_1032 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [15:0] inflight_1; // @[Monitor.scala 723:35]
  reg [63:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [63:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [63:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93]
  wire [63:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[63:1]}; // @[Monitor.scala 747:146]
  wire  _T_1058 = io_in_d_valid & d_first_2 & _T_770; // @[Monitor.scala 779:71]
  wire [15:0] d_clr_1 = _d_first_T & d_first_2 & _T_770 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [142:0] _GEN_68 = _d_first_T & d_first_2 & _T_770 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire [15:0] _T_1066 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_1076 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [15:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [15:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [63:0] d_opcodes_clr_1 = _GEN_68[63:0];
  wire [63:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [63:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_1096 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 16'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 64'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 64'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 16'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 64'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_105 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_105 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_163 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_163 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_105 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_105 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_163 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_163 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_367 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_367 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_532 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_532 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_595 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_595 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_595 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_595 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_766 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_766 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_786 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_786 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(sink_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(sink_ok | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_801 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_805 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(sink_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(sink_ok | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_801 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_805 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_838 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_838 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_838 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_838 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_913 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_913 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_921 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_921 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_925 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_925 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_929 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_929 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_937 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_937 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_941 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_941 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_945 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_945 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_949 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_949 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_953 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_953 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_957 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_957 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_966 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_966 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~(_T_989 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~(_T_989 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_995 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_995 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_999 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_999 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1007 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1007 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1011 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1011 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1021 & ~(_T_1023 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1021 & ~(_T_1023 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1032 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1032 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1058 & ~(_T_1066[0] | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1058 & ~(_T_1066[0] | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1058 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1058 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1096 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:102:11)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1096 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  source = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  address = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  d_first_counter = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  opcode_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  param_1 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  sink = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight = _RAND_12[15:0];
  _RAND_13 = {2{`RANDOM}};
  inflight_opcodes = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_sizes = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  watchdog = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  inflight_1 = _RAND_18[15:0];
  _RAND_19 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  watchdog_1 = _RAND_21[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar_1(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [3:0]  auto_in_a_bits_mask,
  input  [31:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output [5:0]  auto_in_d_bits_sink,
  output        auto_in_d_bits_denied,
  output [31:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_1_a_ready,
  output        auto_out_1_a_valid,
  output [2:0]  auto_out_1_a_bits_opcode,
  output [2:0]  auto_out_1_a_bits_size,
  output [3:0]  auto_out_1_a_bits_source,
  output [12:0] auto_out_1_a_bits_address,
  output [3:0]  auto_out_1_a_bits_mask,
  output        auto_out_1_d_ready,
  input         auto_out_1_d_valid,
  input  [2:0]  auto_out_1_d_bits_opcode,
  input  [2:0]  auto_out_1_d_bits_size,
  input  [3:0]  auto_out_1_d_bits_source,
  input         auto_out_1_d_bits_denied,
  input         auto_out_1_d_bits_corrupt,
  input         auto_out_0_a_ready,
  output        auto_out_0_a_valid,
  output [2:0]  auto_out_0_a_bits_opcode,
  output [2:0]  auto_out_0_a_bits_size,
  output [3:0]  auto_out_0_a_bits_source,
  output [31:0] auto_out_0_a_bits_address,
  output [3:0]  auto_out_0_a_bits_mask,
  output [31:0] auto_out_0_a_bits_data,
  output        auto_out_0_d_ready,
  input         auto_out_0_d_valid,
  input  [2:0]  auto_out_0_d_bits_opcode,
  input  [1:0]  auto_out_0_d_bits_param,
  input  [2:0]  auto_out_0_d_bits_size,
  input  [3:0]  auto_out_0_d_bits_source,
  input  [4:0]  auto_out_0_d_bits_sink,
  input         auto_out_0_d_bits_denied,
  input  [31:0] auto_out_0_d_bits_data,
  input         auto_out_0_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  reg [3:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 4'h0; // @[Arbiter.scala 88:28]
  wire [1:0] readys_filter_lo = {auto_out_1_d_valid,auto_out_0_d_valid}; // @[Cat.scala 30:58]
  reg [1:0] readys_mask; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 24:30]
  wire [1:0] readys_filter_hi = readys_filter_lo & _readys_filter_T; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter = {readys_filter_hi,auto_out_1_d_valid,auto_out_0_d_valid}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_1 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_1; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_2 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready = _GEN_2 | _readys_unready_T_4; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  wire  readys_0 = readys_readys[0]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_0 = readys_0 & auto_out_0_d_valid; // @[Arbiter.scala 97:79]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire [3:0] _T_36 = muxStateEarly_0 ? auto_out_0_d_bits_source : 4'h0; // @[Mux.scala 27:72]
  wire  readys_1 = readys_readys[1]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_1 = readys_1 & auto_out_1_d_valid; // @[Arbiter.scala 97:79]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire [3:0] _T_37 = muxStateEarly_1 ? auto_out_1_d_bits_source : 4'h0; // @[Mux.scala 27:72]
  wire [31:0] _requestAIO_T = auto_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_1 = {1'b0,$signed(_requestAIO_T)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_3 = $signed(_requestAIO_T_1) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_4 = $signed(_requestAIO_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_5 = auto_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_6 = {1'b0,$signed(_requestAIO_T_5)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_8 = $signed(_requestAIO_T_6) & 33'she0000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_9 = $signed(_requestAIO_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_10 = auto_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_11 = {1'b0,$signed(_requestAIO_T_10)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_13 = $signed(_requestAIO_T_11) & 33'shc0000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_14 = $signed(_requestAIO_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_15 = auto_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_16 = {1'b0,$signed(_requestAIO_T_15)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_18 = $signed(_requestAIO_T_16) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  _requestAIO_T_19 = $signed(_requestAIO_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  wire  requestAIO_0_0 = _requestAIO_T_4 | _requestAIO_T_9 | _requestAIO_T_14 | _requestAIO_T_19; // @[Xbar.scala 363:92]
  wire [32:0] _requestAIO_T_24 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_26 = $signed(_requestAIO_T_24) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_1 = $signed(_requestAIO_T_26) == 33'sh0; // @[Parameters.scala 137:67]
  wire [12:0] _beatsDO_decode_T_1 = 13'h3f << auto_out_0_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_3 = ~_beatsDO_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] beatsDO_decode = _beatsDO_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata = auto_out_0_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [3:0] beatsDO_0 = beatsDO_opdata ? beatsDO_decode : 4'h0; // @[Edges.scala 220:14]
  wire [12:0] _beatsDO_decode_T_5 = 13'h3f << auto_out_1_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_7 = ~_beatsDO_decode_T_5[5:0]; // @[package.scala 234:46]
  wire [3:0] beatsDO_decode_1 = _beatsDO_decode_T_7[5:2]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata_1 = auto_out_1_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [3:0] beatsDO_1 = beatsDO_opdata_1 ? beatsDO_decode_1 : 4'h0; // @[Edges.scala 220:14]
  wire  latch = idle & auto_in_d_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _readys_mask_T = readys_readys & readys_filter_lo; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 244:43]
  wire  _prefixOR_T = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 104:53]
  wire  _T_10 = auto_out_0_d_valid | auto_out_1_d_valid; // @[Arbiter.scala 107:36]
  wire  _T_11 = ~(auto_out_0_d_valid | auto_out_1_d_valid); // @[Arbiter.scala 107:15]
  wire [3:0] maskedBeats_0 = earlyWinner_0 ? beatsDO_0 : 4'h0; // @[Arbiter.scala 111:73]
  wire [3:0] maskedBeats_1 = earlyWinner_1 ? beatsDO_1 : 4'h0; // @[Arbiter.scala 111:73]
  wire [3:0] initBeats = maskedBeats_0 | maskedBeats_1; // @[Arbiter.scala 112:44]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & auto_out_0_d_valid | state_1 & auto_out_1_d_valid; // @[Mux.scala 27:72]
  wire  sink_ACancel_5_earlyValid = idle ? _T_10 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_5_earlyValid; // @[ReadyValidCancel.scala 50:33]
  wire [3:0] _GEN_3 = {{3'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [3:0] _beatsLeft_T_4 = beatsLeft - _GEN_3; // @[Arbiter.scala 113:52]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire [5:0] out_1_0_d_bits_sink = {{1'd0}, auto_out_0_d_bits_sink}; // @[Xbar.scala 288:19 Xbar.scala 323:28]
  wire [5:0] _T_33 = muxStateEarly_0 ? out_1_0_d_bits_sink : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_34 = muxStateEarly_1 ? 6'h20 : 6'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_39 = muxStateEarly_0 ? auto_out_0_d_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_40 = muxStateEarly_1 ? auto_out_1_d_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_45 = muxStateEarly_0 ? auto_out_0_d_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_46 = muxStateEarly_1 ? auto_out_1_d_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  TLMonitor_1 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  assign auto_in_a_ready = requestAIO_0_0 & auto_out_0_a_ready | requestAIO_0_1 & auto_out_1_a_ready; // @[Mux.scala 27:72]
  assign auto_in_d_valid = idle ? _T_10 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_in_d_bits_opcode = _T_45 | _T_46; // @[Mux.scala 27:72]
  assign auto_in_d_bits_param = muxStateEarly_0 ? auto_out_0_d_bits_param : 2'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_size = _T_39 | _T_40; // @[Mux.scala 27:72]
  assign auto_in_d_bits_source = _T_36 | _T_37; // @[Mux.scala 27:72]
  assign auto_in_d_bits_sink = _T_33 | _T_34; // @[Mux.scala 27:72]
  assign auto_in_d_bits_denied = muxStateEarly_0 & auto_out_0_d_bits_denied | muxStateEarly_1 & auto_out_1_d_bits_denied
    ; // @[Mux.scala 27:72]
  assign auto_in_d_bits_data = muxStateEarly_0 ? auto_out_0_d_bits_data : 32'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_corrupt = muxStateEarly_0 & auto_out_0_d_bits_corrupt | muxStateEarly_1 &
    auto_out_1_d_bits_corrupt; // @[Mux.scala 27:72]
  assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1; // @[Xbar.scala 428:50]
  assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_1_a_bits_address = auto_in_a_bits_address[12:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_1_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_d_ready = auto_in_d_ready & allowed_1; // @[Arbiter.scala 123:31]
  assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0; // @[Xbar.scala 428:50]
  assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_0_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_d_ready = auto_in_d_ready & allowed_0; // @[Arbiter.scala 123:31]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = requestAIO_0_0 & auto_out_0_a_ready | requestAIO_0_1 & auto_out_1_a_ready; // @[Mux.scala 27:72]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = idle ? _T_10 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign monitor_io_in_d_bits_opcode = _T_45 | _T_46; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_param = muxStateEarly_0 ? auto_out_0_d_bits_param : 2'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_size = _T_39 | _T_40; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_source = _T_36 | _T_37; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_sink = _T_33 | _T_34; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_denied = muxStateEarly_0 & auto_out_0_d_bits_denied | muxStateEarly_1 &
    auto_out_1_d_bits_denied; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_corrupt = muxStateEarly_0 & auto_out_0_d_bits_corrupt | muxStateEarly_1 &
    auto_out_1_d_bits_corrupt; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 4'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin // @[Arbiter.scala 113:23]
      beatsLeft <= initBeats;
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch & |readys_filter_lo) begin // @[Arbiter.scala 27:32]
      readys_mask <= _readys_mask_T_3; // @[Arbiter.scala 28:12]
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin // @[Arbiter.scala 117:30]
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin // @[Arbiter.scala 117:30]
      state_1 <= earlyWinner_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(auto_out_0_d_valid | auto_out_1_d_valid) | _prefixOR_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(auto_out_0_d_valid | auto_out_1_d_valid) | _prefixOR_T | reset)) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_11 | _T_10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_11 | _T_10 | reset)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  readys_mask = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  state_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_2(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [3:0]  io_in_a_bits_source,
  input  [12:0] io_in_a_bits_address,
  input  [3:0]  io_in_a_bits_mask,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [2:0]  io_in_d_bits_size,
  input  [3:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = ~io_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | io_in_a_bits_source[3]; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [12:0] _GEN_71 = {{7'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [12:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 13'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_34 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_54 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [12:0] _T_57 = io_in_a_bits_address ^ 13'h1000; // @[Parameters.scala 137:31]
  wire [13:0] _T_58 = {1'b0,$signed(_T_57)}; // @[Parameters.scala 137:49]
  wire [13:0] _T_60 = $signed(_T_58) & -14'sh1000; // @[Parameters.scala 137:52]
  wire  _T_61 = $signed(_T_60) == 14'sh0; // @[Parameters.scala 137:67]
  wire  _T_62 = _T_54 & _T_61; // @[Parameters.scala 670:56]
  wire  _T_64 = source_ok & _T_62; // @[Monitor.scala 82:72]
  wire [3:0] _T_97 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_98 = _T_97 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_106 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_182 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_228 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_236 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_284 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_328 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_329 = io_in_a_bits_mask & _T_328; // @[Monitor.scala 127:31]
  wire  _T_330 = _T_329 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_334 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_382 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_430 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_482 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_13 = ~io_in_d_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_13 | io_in_d_bits_source[3]; // @[Parameters.scala 1125:46]
  wire  _T_486 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_490 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_498 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_502 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_506 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_534 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_554 = _T_502 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_563 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_580 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_598 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [3:0] source; // @[Monitor.scala 387:22]
  reg [12:0] address; // @[Monitor.scala 388:22]
  wire  _T_628 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_629 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_637 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_641 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_645 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [3:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_652 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_653 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_661 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_665 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_673 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [15:0] inflight; // @[Monitor.scala 611:27]
  reg [63:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [63:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69]
  wire [63:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [63:0] _GEN_73 = {{48'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[63:1]}; // @[Monitor.scala 634:152]
  wire [63:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [63:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91]
  wire [63:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[63:1]}; // @[Monitor.scala 638:144]
  wire  _T_679 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [15:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_682 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [15:0] _T_684 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_686 = ~_T_684[0]; // @[Monitor.scala 658:17]
  wire [15:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [130:0] _GEN_19 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [130:0] _GEN_20 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_690 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_692 = ~_T_486; // @[Monitor.scala 671:74]
  wire  _T_693 = io_in_d_valid & d_first_1 & ~_T_486; // @[Monitor.scala 671:71]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [15:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_486 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [15:0] d_clr = _d_first_T & d_first_1 & _T_692 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [142:0] _GEN_23 = _d_first_T & d_first_1 & _T_692 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_679 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [15:0] _T_703 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_705 = _T_703[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_710 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39]
  wire  _T_711 = io_in_d_bits_opcode == _GEN_32 | _T_710; // @[Monitor.scala 685:77]
  wire  _T_715 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_722 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_723 = io_in_d_bits_opcode == _GEN_48 | _T_722; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_727 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_737 = _T_690 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_692; // @[Monitor.scala 694:116]
  wire  _T_739 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_746 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [15:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [15:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [15:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [63:0] a_opcodes_set = _GEN_19[63:0];
  wire [63:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [63:0] d_opcodes_clr = _GEN_23[63:0];
  wire [63:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [63:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [63:0] a_sizes_set = _GEN_20[63:0];
  wire [63:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [63:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_755 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [15:0] inflight_1; // @[Monitor.scala 723:35]
  reg [63:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [63:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [63:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93]
  wire [63:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[63:1]}; // @[Monitor.scala 747:146]
  wire  _T_781 = io_in_d_valid & d_first_2 & _T_486; // @[Monitor.scala 779:71]
  wire [15:0] d_clr_1 = _d_first_T & d_first_2 & _T_486 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [142:0] _GEN_68 = _d_first_T & d_first_2 & _T_486 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire [15:0] _T_789 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_799 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [15:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [15:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [63:0] d_opcodes_clr_1 = _GEN_68[63:0];
  wire [63:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [63:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_824 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 16'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 64'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 64'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 16'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 64'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_98 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_98 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_T_98 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_T_98 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_62 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_62 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(_T_330 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(_T_330 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_482 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_482 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_490 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_490 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_498 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_498 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_502 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_502 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(_T_490 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(_T_490 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(_T_498 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(_T_498 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(_T_490 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(_T_490 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(_T_554 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(_T_554 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_563 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_563 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_563 & ~(_T_498 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_563 & ~(_T_498 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_580 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_580 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_580 & ~(_T_554 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_580 & ~(_T_554 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_598 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_598 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_598 & ~(_T_498 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_598 & ~(_T_498 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628 & ~(_T_629 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628 & ~(_T_629 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628 & ~(_T_637 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628 & ~(_T_637 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628 & ~(_T_641 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628 & ~(_T_641 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628 & ~(_T_645 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628 & ~(_T_645 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & ~(_T_653 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & ~(_T_653 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & ~(_T_661 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & ~(_T_661 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & ~(_T_665 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & ~(_T_665 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & ~(_T_673 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & ~(_T_673 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_682 & ~(_T_686 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_682 & ~(_T_686 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & ~(_T_705 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & ~(_T_705 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & same_cycle_resp & ~(_T_711 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & same_cycle_resp & ~(_T_711 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & same_cycle_resp & ~(_T_715 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & same_cycle_resp & ~(_T_715 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & ~same_cycle_resp & ~(_T_723 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & ~same_cycle_resp & ~(_T_723 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & ~same_cycle_resp & ~(_T_727 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & ~same_cycle_resp & ~(_T_727 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_737 & ~(_T_739 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_737 & ~(_T_739 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_746 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_746 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_755 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_755 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_781 & ~(_T_789[0] | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_781 & ~(_T_789[0] | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_781 & ~(_T_799 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_781 & ~(_T_799 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_824 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:43:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_824 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  source = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  address = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  d_first_counter = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  opcode_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  size_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  source_1 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  denied = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  inflight = _RAND_10[15:0];
  _RAND_11 = {2{`RANDOM}};
  inflight_opcodes = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  inflight_sizes = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  watchdog = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  inflight_1 = _RAND_16[15:0];
  _RAND_17 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  watchdog_1 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [2:0] io_enq_bits_size,
  input  [3:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_size,
  output [3:0] io_deq_bits_source
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] ram_source [0:0]; // @[Decoupled.scala 218:16]
  wire [3:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign ram_opcode_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = 1'h0;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = 1'h0;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLError(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [12:0] auto_in_a_bits_address,
  input  [3:0]  auto_in_a_bits_mask,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output        auto_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [12:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  a_clock; // @[Decoupled.scala 296:21]
  wire  a_reset; // @[Decoupled.scala 296:21]
  wire  a_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  a_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] a_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] a_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [3:0] a_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire  a_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  a_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] a_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] a_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [3:0] a_io_deq_bits_source; // @[Decoupled.scala 296:21]
  reg  idle; // @[Error.scala 44:23]
  wire  _a_last_T = a_io_deq_ready & a_io_deq_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _a_last_beats1_decode_T_1 = 13'h3f << a_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] _a_last_beats1_decode_T_3 = ~_a_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] a_last_beats1_decode = _a_last_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  a_last_beats1_opdata = ~a_io_deq_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [3:0] a_last_beats1 = a_last_beats1_opdata ? a_last_beats1_decode : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] a_last_counter; // @[Edges.scala 228:27]
  wire [3:0] a_last_counter1 = a_last_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_last_first = a_last_counter == 4'h0; // @[Edges.scala 230:25]
  wire  a_last = a_last_counter == 4'h1 | a_last_beats1 == 4'h0; // @[Edges.scala 231:37]
  reg [3:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle_1 = beatsLeft == 4'h0; // @[Arbiter.scala 88:28]
  wire  da_valid = a_io_deq_valid & a_last & idle; // @[Error.scala 51:35]
  wire [1:0] _readys_T = {da_valid,1'h0}; // @[Cat.scala 30:58]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[package.scala 244:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[Arbiter.scala 16:61]
  wire  readys_1 = _readys_T_7[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle_1 ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_in_d_ready & allowed_1; // @[Arbiter.scala 123:31]
  wire  _T = out_1_ready & da_valid; // @[Decoupled.scala 40:37]
  wire [2:0] da_bits_size = a_io_deq_bits_size; // @[Error.scala 43:18 Error.scala 55:21]
  wire [12:0] _beats1_decode_T_1 = 13'h3f << da_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] beats1_decode = _beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire [2:0] _GEN_4 = 3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_5 = 3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_4; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_6 = 3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_5; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_7 = 3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_6; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_8 = 3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_7; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] da_bits_opcode = 3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8; // @[Error.scala 53:21 Error.scala 53:21]
  wire  beats1_opdata = da_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [3:0] beats1 = beats1_opdata ? beats1_decode : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] counter; // @[Edges.scala 228:27]
  wire [3:0] counter1 = counter - 4'h1; // @[Edges.scala 229:28]
  wire  da_first = counter == 4'h0; // @[Edges.scala 230:25]
  wire  da_last = counter == 4'h1 | beats1 == 4'h0; // @[Edges.scala 231:37]
  wire  _GEN_12 = _T & da_bits_opcode == 3'h4 ? 1'h0 : idle; // @[Error.scala 70:52 Error.scala 70:59 Error.scala 44:23]
  wire  latch = idle_1 & auto_in_d_ready; // @[Arbiter.scala 89:24]
  wire  earlyWinner_1 = readys_1 & da_valid; // @[Arbiter.scala 97:79]
  wire  _T_22 = ~da_valid; // @[Arbiter.scala 107:15]
  wire  muxStateEarly_1 = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_2 = state_1 & da_valid; // @[Mux.scala 27:72]
  wire  sink_ACancel_earlyValid = idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 50:33]
  wire [3:0] _GEN_17 = {{3'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [3:0] _beatsLeft_T_4 = beatsLeft - _GEN_17; // @[Arbiter.scala 113:52]
  wire [3:0] da_bits_source = a_io_deq_bits_source; // @[Error.scala 43:18 Error.scala 56:21]
  TLMonitor_2 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue a ( // @[Decoupled.scala 296:21]
    .clock(a_clock),
    .reset(a_reset),
    .io_enq_ready(a_io_enq_ready),
    .io_enq_valid(a_io_enq_valid),
    .io_enq_bits_opcode(a_io_enq_bits_opcode),
    .io_enq_bits_size(a_io_enq_bits_size),
    .io_enq_bits_source(a_io_enq_bits_source),
    .io_deq_ready(a_io_deq_ready),
    .io_deq_valid(a_io_deq_valid),
    .io_deq_bits_opcode(a_io_deq_bits_opcode),
    .io_deq_bits_size(a_io_deq_bits_size),
    .io_deq_bits_source(a_io_deq_bits_source)
  );
  assign auto_in_a_ready = a_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign auto_in_d_valid = idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2; // @[Arbiter.scala 125:29]
  assign auto_in_d_bits_opcode = muxStateEarly_1 ? da_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_size = muxStateEarly_1 ? da_bits_size : 3'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_source = muxStateEarly_1 ? da_bits_source : 4'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_denied = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  assign auto_in_d_bits_corrupt = muxStateEarly_1 & beats1_opdata; // @[Mux.scala 27:72]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = a_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2; // @[Arbiter.scala 125:29]
  assign monitor_io_in_d_bits_opcode = muxStateEarly_1 ? da_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_size = muxStateEarly_1 ? da_bits_size : 3'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_source = muxStateEarly_1 ? da_bits_source : 4'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_denied = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  assign monitor_io_in_d_bits_corrupt = muxStateEarly_1 & beats1_opdata; // @[Mux.scala 27:72]
  assign a_clock = clock;
  assign a_reset = reset;
  assign a_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_deq_ready = out_1_ready & da_last & idle | ~a_last; // @[Error.scala 50:46]
  always @(posedge clock) begin
    idle <= reset | _GEN_12; // @[Error.scala 44:23 Error.scala 44:23]
    if (reset) begin // @[Edges.scala 228:27]
      a_last_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_last_T) begin // @[Edges.scala 234:17]
      if (a_last_first) begin // @[Edges.scala 235:21]
        if (a_last_beats1_opdata) begin // @[Edges.scala 220:14]
          a_last_counter <= a_last_beats1_decode;
        end else begin
          a_last_counter <= 4'h0;
        end
      end else begin
        a_last_counter <= a_last_counter1;
      end
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 4'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin // @[Arbiter.scala 113:23]
      if (earlyWinner_1) begin // @[Arbiter.scala 111:73]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          beatsLeft <= beats1_decode;
        end else begin
          beatsLeft <= 4'h0;
        end
      end else begin
        beatsLeft <= 4'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin // @[Arbiter.scala 117:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T) begin // @[Edges.scala 234:17]
      if (da_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          counter <= beats1_decode;
        end else begin
          counter <= 4'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(idle | da_first | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Error.scala:49 assert (idle || da_first) // we only send Grant, never GrantData => simplified flow control below\n"
            ); // @[Error.scala 49:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(idle | da_first | reset)) begin
          $fatal; // @[Error.scala 49:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~da_valid | earlyWinner_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~da_valid | earlyWinner_1 | reset)) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_22 | da_valid | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_22 | da_valid | reset)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  idle = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  a_last_counter = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  beatsLeft = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  state_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  counter = _RAND_4[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_3(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [3:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [3:0]  io_in_a_bits_mask,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [3:0]  io_in_d_bits_source,
  input  [4:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = ~io_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | io_in_a_bits_source[3]; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_34 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_60 = 3'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48]
  wire [31:0] _T_62 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_63 = {1'b0,$signed(_T_62)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_65 = $signed(_T_63) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_66 = $signed(_T_65) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_77 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_78 = {1'b0,$signed(_T_77)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_80 = $signed(_T_78) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_81 = $signed(_T_80) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_82 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_83 = {1'b0,$signed(_T_82)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_85 = $signed(_T_83) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_86 = $signed(_T_85) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_90 = _T_66 | _T_71 | _T_76 | _T_81 | _T_86; // @[Parameters.scala 671:42]
  wire  _T_91 = _T_60 & _T_90; // @[Parameters.scala 670:56]
  wire  _T_94 = source_ok & _T_91; // @[Monitor.scala 82:72]
  wire [32:0] _T_120 = $signed(_T_78) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _T_121 = $signed(_T_120) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_124 = _T_66 | _T_71 | _T_76 | _T_121; // @[Parameters.scala 671:42]
  wire [3:0] _T_145 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_146 = _T_145 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_154 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_278 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_301 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_327 = _T_301 & _T_124; // @[Parameters.scala 670:56]
  wire  _T_342 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_350 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_398 = source_ok & _T_327; // @[Monitor.scala 115:71]
  wire  _T_416 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_478 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_479 = io_in_a_bits_mask & _T_478; // @[Monitor.scala 127:31]
  wire  _T_480 = _T_479 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_484 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_504 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_530 = _T_504 & _T_124; // @[Parameters.scala 670:56]
  wire  _T_532 = source_ok & _T_530; // @[Monitor.scala 131:74]
  wire  _T_550 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_616 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_686 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_13 = ~io_in_d_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_13 | io_in_d_bits_source[3]; // @[Parameters.scala 1125:46]
  wire  _T_690 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_694 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_698 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_702 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_706 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_710 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_721 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_725 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_738 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_758 = _T_706 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_767 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_784 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_802 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [3:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_832 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_833 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_841 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_845 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_849 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [3:0] source_1; // @[Monitor.scala 538:22]
  reg [4:0] sink; // @[Monitor.scala 539:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_856 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_857 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_861 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_865 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_869 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_873 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29]
  wire  _T_877 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [15:0] inflight; // @[Monitor.scala 611:27]
  reg [63:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [63:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69]
  wire [63:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [63:0] _GEN_73 = {{48'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[63:1]}; // @[Monitor.scala 634:152]
  wire [63:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [63:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91]
  wire [63:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[63:1]}; // @[Monitor.scala 638:144]
  wire  _T_883 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire  _T_886 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [15:0] _T_888 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_890 = ~_T_888[0]; // @[Monitor.scala 658:17]
  wire [15:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [130:0] _GEN_19 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [130:0] _GEN_20 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_894 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_896 = ~_T_690; // @[Monitor.scala 671:74]
  wire  _T_897 = io_in_d_valid & d_first_1 & ~_T_690; // @[Monitor.scala 671:71]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [15:0] d_clr = _d_first_T & d_first_1 & _T_896 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [142:0] _GEN_23 = _d_first_T & d_first_1 & _T_896 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_883 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [15:0] _T_907 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_909 = _T_907[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_914 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39]
  wire  _T_915 = io_in_d_bits_opcode == _GEN_32 | _T_914; // @[Monitor.scala 685:77]
  wire  _T_919 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_926 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_927 = io_in_d_bits_opcode == _GEN_48 | _T_926; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_931 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_941 = _T_894 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_896; // @[Monitor.scala 694:116]
  wire  _T_943 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire [15:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [15:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [15:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [63:0] a_opcodes_set = _GEN_19[63:0];
  wire [63:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [63:0] d_opcodes_clr = _GEN_23[63:0];
  wire [63:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [63:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [63:0] a_sizes_set = _GEN_20[63:0];
  wire [63:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [63:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_952 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [15:0] inflight_1; // @[Monitor.scala 723:35]
  reg [63:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [63:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [63:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93]
  wire [63:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[63:1]}; // @[Monitor.scala 747:146]
  wire  _T_978 = io_in_d_valid & d_first_2 & _T_690; // @[Monitor.scala 779:71]
  wire [15:0] d_clr_1 = _d_first_T & d_first_2 & _T_690 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [142:0] _GEN_68 = _d_first_T & d_first_2 & _T_690 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire [15:0] _T_986 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_996 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [15:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [15:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [63:0] d_opcodes_clr_1 = _GEN_68[63:0];
  wire [63:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [63:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_1016 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 16'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 64'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 64'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 16'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 64'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_94 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_94 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_146 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_146 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_T_94 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_T_94 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_T_146 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_T_146 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(_T_327 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(_T_327 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(_T_398 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(_T_398 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(_T_398 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(_T_398 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(_T_480 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(_T_480 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(_T_532 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(_T_532 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(_T_532 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(_T_532 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(_T_398 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(_T_398 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_686 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_686 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_694 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_694 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_698 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_698 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_702 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_702 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_706 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_706 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_694 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_694 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_721 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_725 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_725 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_702 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_702 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_694 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_694 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_721 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_725 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_725 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_758 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_758 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(_T_698 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(_T_698 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(_T_702 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(_T_702 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(_T_698 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(_T_698 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(_T_758 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(_T_758 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(_T_698 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(_T_698 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(_T_702 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(_T_702 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & ~(_T_833 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & ~(_T_833 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & ~(_T_841 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & ~(_T_841 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & ~(_T_845 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & ~(_T_845 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & ~(_T_849 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & ~(_T_849 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_857 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_857 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_861 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_861 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_865 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_865 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_869 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_869 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_873 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_873 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_877 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_877 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_886 & ~(_T_890 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_886 & ~(_T_890 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & ~(_T_909 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & ~(_T_909 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & same_cycle_resp & ~(_T_915 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & same_cycle_resp & ~(_T_915 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & same_cycle_resp & ~(_T_919 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & same_cycle_resp & ~(_T_919 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & ~same_cycle_resp & ~(_T_927 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & ~same_cycle_resp & ~(_T_927 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & ~same_cycle_resp & ~(_T_931 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & ~same_cycle_resp & ~(_T_931 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_941 & ~(_T_943 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_941 & ~(_T_943 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_952 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_952 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_978 & ~(_T_986[0] | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_978 & ~(_T_986[0] | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_978 & ~(_T_996 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_978 & ~(_T_996 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1016 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1016 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  source = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  address = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  d_first_counter = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  opcode_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  param_1 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  sink = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight = _RAND_12[15:0];
  _RAND_13 = {2{`RANDOM}};
  inflight_opcodes = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_sizes = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  watchdog = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  inflight_1 = _RAND_18[15:0];
  _RAND_19 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  watchdog_1 = _RAND_21[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBusBypassBar(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [2:0]   auto_in_a_bits_size,
  input  [3:0]   auto_in_a_bits_source,
  input  [31:0]  auto_in_a_bits_address,
  input  [3:0]   auto_in_a_bits_mask,
  input  [31:0]  auto_in_a_bits_data,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [2:0]   auto_in_d_bits_opcode,
  output [1:0]   auto_in_d_bits_param,
  output [2:0]   auto_in_d_bits_size,
  output [3:0]   auto_in_d_bits_source,
  output [4:0]   auto_in_d_bits_sink,
  output         auto_in_d_bits_denied,
  output [31:0]  auto_in_d_bits_data,
  output         auto_in_d_bits_corrupt,
  input          auto_out_1_a_ready,
  output         auto_out_1_a_valid,
  output [2:0]   auto_out_1_a_bits_opcode,
  output [2:0]   auto_out_1_a_bits_size,
  output [3:0]   auto_out_1_a_bits_source,
  output [31:0]  auto_out_1_a_bits_address,
  output [3:0]   auto_out_1_a_bits_mask,
  output [31:0]  auto_out_1_a_bits_data,
  output         auto_out_1_d_ready,
  input          auto_out_1_d_valid,
  input  [2:0]   auto_out_1_d_bits_opcode,
  input  [1:0]   auto_out_1_d_bits_param,
  input  [2:0]   auto_out_1_d_bits_size,
  input  [3:0]   auto_out_1_d_bits_source,
  input  [4:0]   auto_out_1_d_bits_sink,
  input          auto_out_1_d_bits_denied,
  input  [31:0]  auto_out_1_d_bits_data,
  input          auto_out_1_d_bits_corrupt,
  input          auto_out_0_a_ready,
  output         auto_out_0_a_valid,
  output [2:0]   auto_out_0_a_bits_opcode,
  output [3:0]   auto_out_0_a_bits_size,
  output [3:0]   auto_out_0_a_bits_source,
  output [127:0] auto_out_0_a_bits_address,
  output [3:0]   auto_out_0_a_bits_mask,
  output         auto_out_0_d_ready,
  input          auto_out_0_d_valid,
  input  [2:0]   auto_out_0_d_bits_opcode,
  input  [3:0]   auto_out_0_d_bits_size,
  input  [3:0]   auto_out_0_d_bits_source,
  input          auto_out_0_d_bits_denied,
  input          auto_out_0_d_bits_corrupt,
  input          io_bypass
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire [4:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  reg  in_reset; // @[BusBypass.scala 77:27]
  reg  bypass_reg; // @[BusBypass.scala 78:25]
  wire  bypass = in_reset ? io_bypass : bypass_reg; // @[BusBypass.scala 79:21]
  reg [5:0] flight; // @[Edges.scala 294:25]
  reg [3:0] stall_counter; // @[Edges.scala 228:27]
  wire  stall_first = stall_counter == 4'h0; // @[Edges.scala 230:25]
  wire  stall = bypass != io_bypass & stall_first; // @[BusBypass.scala 84:40]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[BusBypass.scala 88:21]
  wire  _bundleIn_0_a_ready_T_1 = bypass ? auto_out_0_a_ready : auto_out_1_a_ready; // @[BusBypass.scala 88:34]
  wire  in_a_ready = ~stall & _bundleIn_0_a_ready_T_1; // @[BusBypass.scala 88:28]
  wire  _T = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _beats1_decode_T_1 = 13'h3f << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] beats1_decode = _beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] counter; // @[Edges.scala 228:27]
  wire [3:0] counter1 = counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = counter == 4'h0; // @[Edges.scala 230:25]
  wire  in_d_valid = bypass ? auto_out_0_d_valid : auto_out_1_d_valid; // @[BusBypass.scala 94:24]
  wire  _T_3 = auto_in_d_ready & in_d_valid; // @[Decoupled.scala 40:37]
  wire [2:0] bundleIn_0_d_bits_out_size = auto_out_0_d_bits_size[2:0]; // @[BusBypass.scala 95:46 BusBypass.scala 95:63]
  wire [2:0] in_d_bits_size = bypass ? bundleIn_0_d_bits_out_size : auto_out_1_d_bits_size; // @[BusBypass.scala 96:21]
  wire [12:0] _beats1_decode_T_13 = 13'h3f << in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_15 = ~_beats1_decode_T_13[5:0]; // @[package.scala 234:46]
  wire [3:0] beats1_decode_3 = _beats1_decode_T_15[5:2]; // @[Edges.scala 219:59]
  wire [2:0] in_d_bits_opcode = bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode; // @[BusBypass.scala 96:21]
  wire  beats1_opdata_3 = in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [3:0] beats1_3 = beats1_opdata_3 ? beats1_decode_3 : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] counter_3; // @[Edges.scala 228:27]
  wire [3:0] counter1_3 = counter_3 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = counter_3 == 4'h0; // @[Edges.scala 230:25]
  wire  d_last = counter_3 == 4'h1 | beats1_3 == 4'h0; // @[Edges.scala 231:37]
  wire  d_request = in_d_bits_opcode[2] & ~in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  inc_hi = _T & a_first; // @[Edges.scala 309:28]
  wire  inc_lo = _T_3 & d_first & d_request; // @[Edges.scala 312:39]
  wire [1:0] inc = {inc_hi,inc_lo}; // @[Cat.scala 30:58]
  wire  dec_lo = _T_3 & d_last; // @[Edges.scala 319:28]
  wire [1:0] dec = {1'h0,dec_lo}; // @[Cat.scala 30:58]
  wire [1:0] _next_flight_T_2 = inc[0] + inc[1]; // @[Bitwise.scala 47:55]
  wire [5:0] _GEN_7 = {{4'd0}, _next_flight_T_2}; // @[Edges.scala 323:30]
  wire [5:0] _next_flight_T_5 = flight + _GEN_7; // @[Edges.scala 323:30]
  wire [1:0] _next_flight_T_8 = dec[0] + dec[1]; // @[Bitwise.scala 47:55]
  wire [5:0] _GEN_8 = {{4'd0}, _next_flight_T_8}; // @[Edges.scala 323:46]
  wire [5:0] next_flight = _next_flight_T_5 - _GEN_8; // @[Edges.scala 323:46]
  wire [3:0] stall_counter1 = stall_counter - 4'h1; // @[Edges.scala 229:28]
  wire  _bundleOut_0_a_valid_T_1 = _bundleIn_0_a_ready_T & auto_in_a_valid; // @[BusBypass.scala 86:28]
  wire  _bundleOut_1_a_valid_T_2 = ~bypass; // @[BusBypass.scala 87:45]
  TLMonitor_3 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  assign auto_in_a_ready = ~stall & _bundleIn_0_a_ready_T_1; // @[BusBypass.scala 88:28]
  assign auto_in_d_valid = bypass ? auto_out_0_d_valid : auto_out_1_d_valid; // @[BusBypass.scala 94:24]
  assign auto_in_d_bits_opcode = bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode; // @[BusBypass.scala 96:21]
  assign auto_in_d_bits_param = bypass ? 2'h0 : auto_out_1_d_bits_param; // @[BusBypass.scala 96:21]
  assign auto_in_d_bits_size = bypass ? bundleIn_0_d_bits_out_size : auto_out_1_d_bits_size; // @[BusBypass.scala 96:21]
  assign auto_in_d_bits_source = bypass ? auto_out_0_d_bits_source : auto_out_1_d_bits_source; // @[BusBypass.scala 96:21]
  assign auto_in_d_bits_sink = bypass ? 5'h0 : auto_out_1_d_bits_sink; // @[BusBypass.scala 96:21]
  assign auto_in_d_bits_denied = bypass ? auto_out_0_d_bits_denied : auto_out_1_d_bits_denied; // @[BusBypass.scala 96:21]
  assign auto_in_d_bits_data = bypass ? 32'h0 : auto_out_1_d_bits_data; // @[BusBypass.scala 96:21]
  assign auto_in_d_bits_corrupt = bypass ? auto_out_0_d_bits_corrupt : auto_out_1_d_bits_corrupt; // @[BusBypass.scala 96:21]
  assign auto_out_1_a_valid = _bundleOut_0_a_valid_T_1 & ~bypass; // @[BusBypass.scala 87:42]
  assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_d_ready = auto_in_d_ready & _bundleOut_1_a_valid_T_2; // @[BusBypass.scala 93:32]
  assign auto_out_0_a_valid = _bundleIn_0_a_ready_T & auto_in_a_valid & bypass; // @[BusBypass.scala 86:42]
  assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_size = {{1'd0}, auto_in_a_bits_size}; // @[Nodes.scala 1207:84 BusBypass.scala 89:18]
  assign auto_out_0_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_address = {{96'd0}, auto_in_a_bits_address}; // @[Nodes.scala 1207:84 BusBypass.scala 89:18]
  assign auto_out_0_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_d_ready = auto_in_d_ready & bypass; // @[BusBypass.scala 92:32]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = ~stall & _bundleIn_0_a_ready_T_1; // @[BusBypass.scala 88:28]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = bypass ? auto_out_0_d_valid : auto_out_1_d_valid; // @[BusBypass.scala 94:24]
  assign monitor_io_in_d_bits_opcode = bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode; // @[BusBypass.scala 96:21]
  assign monitor_io_in_d_bits_param = bypass ? 2'h0 : auto_out_1_d_bits_param; // @[BusBypass.scala 96:21]
  assign monitor_io_in_d_bits_size = bypass ? bundleIn_0_d_bits_out_size : auto_out_1_d_bits_size; // @[BusBypass.scala 96:21]
  assign monitor_io_in_d_bits_source = bypass ? auto_out_0_d_bits_source : auto_out_1_d_bits_source; // @[BusBypass.scala 96:21]
  assign monitor_io_in_d_bits_sink = bypass ? 5'h0 : auto_out_1_d_bits_sink; // @[BusBypass.scala 96:21]
  assign monitor_io_in_d_bits_denied = bypass ? auto_out_0_d_bits_denied : auto_out_1_d_bits_denied; // @[BusBypass.scala 96:21]
  assign monitor_io_in_d_bits_corrupt = bypass ? auto_out_0_d_bits_corrupt : auto_out_1_d_bits_corrupt; // @[BusBypass.scala 96:21]
  always @(posedge clock) begin
    in_reset <= reset; // @[BusBypass.scala 77:27 BusBypass.scala 77:27 BusBypass.scala 77:27]
    if (in_reset | next_flight == 6'h0) begin // @[BusBypass.scala 83:50]
      bypass_reg <= io_bypass; // @[BusBypass.scala 83:63]
    end
    if (reset) begin // @[Edges.scala 294:25]
      flight <= 6'h0; // @[Edges.scala 294:25]
    end else begin
      flight <= next_flight; // @[Edges.scala 324:12]
    end
    if (reset) begin // @[Edges.scala 228:27]
      stall_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T) begin // @[Edges.scala 234:17]
      if (stall_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          stall_counter <= beats1_decode;
        end else begin
          stall_counter <= 4'h0;
        end
      end else begin
        stall_counter <= stall_counter1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          counter <= beats1_decode;
        end else begin
          counter <= 4'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter_3 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T_3) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata_3) begin // @[Edges.scala 220:14]
          counter_3 <= beats1_decode_3;
        end else begin
          counter_3 <= 4'h0;
        end
      end else begin
        counter_3 <= counter1_3;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_reset = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bypass_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  flight = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  stall_counter = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  counter = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  counter_3 = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_4(
  input          clock,
  input          reset,
  input          io_in_a_ready,
  input          io_in_a_valid,
  input  [2:0]   io_in_a_bits_opcode,
  input  [3:0]   io_in_a_bits_size,
  input  [3:0]   io_in_a_bits_source,
  input  [127:0] io_in_a_bits_address,
  input  [3:0]   io_in_a_bits_mask,
  input          io_in_d_ready,
  input          io_in_d_valid,
  input  [2:0]   io_in_d_bits_opcode,
  input  [3:0]   io_in_d_bits_size,
  input  [3:0]   io_in_d_bits_source,
  input          io_in_d_bits_denied,
  input          io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = ~io_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | io_in_a_bits_source[3]; // @[Parameters.scala 1125:46]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46]
  wire [127:0] _GEN_71 = {{116'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [127:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 128'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 4'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire [128:0] _T_12 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire  _T_34 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_36 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42]
  wire  _T_51 = _T_36 & source_ok; // @[Parameters.scala 1160:30]
  wire [128:0] _T_60 = $signed(_T_12) & 129'sh100000000000000000000000000000000; // @[Parameters.scala 137:52]
  wire  _T_61 = $signed(_T_60) == 129'sh0; // @[Parameters.scala 137:67]
  wire  _T_62 = _T_36 & _T_61; // @[Parameters.scala 670:56]
  wire  _T_64 = _T_51 & _T_62; // @[Monitor.scala 82:72]
  wire [3:0] _T_97 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_98 = _T_97 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_106 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_182 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_228 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_236 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_284 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_328 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_329 = io_in_a_bits_mask & _T_328; // @[Monitor.scala 127:31]
  wire  _T_330 = _T_329 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_334 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_354 = io_in_a_bits_size <= 4'h4; // @[Parameters.scala 92:42]
  wire  _T_362 = _T_354 & _T_61; // @[Parameters.scala 670:56]
  wire  _T_364 = _T_51 & _T_362; // @[Monitor.scala 131:74]
  wire  _T_382 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_430 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_482 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_13 = ~io_in_d_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_13 | io_in_d_bits_source[3]; // @[Parameters.scala 1125:46]
  wire  _T_486 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_490 = io_in_d_bits_size >= 4'h2; // @[Monitor.scala 312:27]
  wire  _T_498 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_502 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_506 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_534 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_554 = _T_502 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_563 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_580 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_598 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [9:0] a_first_counter; // @[Edges.scala 228:27]
  wire [9:0] a_first_counter1 = a_first_counter - 10'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 10'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [3:0] size; // @[Monitor.scala 386:22]
  reg [3:0] source; // @[Monitor.scala 387:22]
  reg [127:0] address; // @[Monitor.scala 388:22]
  wire  _T_628 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_629 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_637 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_641 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_645 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [9:0] d_first_counter; // @[Edges.scala 228:27]
  wire [9:0] d_first_counter1 = d_first_counter - 10'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 10'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [3:0] size_1; // @[Monitor.scala 537:22]
  reg [3:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_652 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_653 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_661 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_665 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_673 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [15:0] inflight; // @[Monitor.scala 611:27]
  reg [63:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [127:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [9:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 10'h0; // @[Edges.scala 230:25]
  reg [9:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 10'h0; // @[Edges.scala 230:25]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69]
  wire [63:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [63:0] _GEN_73 = {{48'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[63:1]}; // @[Monitor.scala 634:152]
  wire [6:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65]
  wire [127:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57]
  wire [127:0] _GEN_75 = {{112'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 638:91]
  wire [127:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_75; // @[Monitor.scala 638:91]
  wire [127:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[127:1]}; // @[Monitor.scala 638:144]
  wire  _T_679 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire  _T_682 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59]
  wire [5:0] _GEN_77 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_77}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [130:0] _GEN_78 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_78 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [6:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 657:77]
  wire [4:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [131:0] _GEN_79 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [131:0] _a_sizes_set_T_1 = _GEN_79 << _a_sizes_set_T; // @[Monitor.scala 657:52]
  wire [15:0] _T_684 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_686 = ~_T_684[0]; // @[Monitor.scala 658:17]
  wire [15:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [130:0] _GEN_19 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [131:0] _GEN_20 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 132'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_690 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_692 = ~_T_486; // @[Monitor.scala 671:74]
  wire  _T_693 = io_in_d_valid & d_first_1 & ~_T_486; // @[Monitor.scala 671:71]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [142:0] _GEN_81 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_81 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [142:0] _GEN_82 = {{127'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74]
  wire [142:0] _d_sizes_clr_T_5 = _GEN_82 << _a_size_lookup_T; // @[Monitor.scala 678:74]
  wire [15:0] d_clr = _d_first_T & d_first_1 & _T_692 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [142:0] _GEN_23 = _d_first_T & d_first_1 & _T_692 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire [142:0] _GEN_24 = _d_first_T & d_first_1 & _T_692 ? _d_sizes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 Monitor.scala 678:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_679 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [15:0] _T_703 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_705 = _T_703[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_710 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39]
  wire  _T_711 = io_in_d_bits_opcode == _GEN_32 | _T_710; // @[Monitor.scala 685:77]
  wire  _T_715 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_722 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_723 = io_in_d_bits_opcode == _GEN_48 | _T_722; // @[Monitor.scala 689:72]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0];
  wire [7:0] _GEN_83 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_727 = _GEN_83 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_737 = _T_690 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_692; // @[Monitor.scala 694:116]
  wire  _T_739 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire [15:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [15:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [15:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [63:0] a_opcodes_set = _GEN_19[63:0];
  wire [63:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [63:0] d_opcodes_clr = _GEN_23[63:0];
  wire [63:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [63:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [127:0] a_sizes_set = _GEN_20[127:0];
  wire [127:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [127:0] d_sizes_clr = _GEN_24[127:0];
  wire [127:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56]
  wire [127:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_748 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [15:0] inflight_1; // @[Monitor.scala 723:35]
  reg [127:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [9:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 10'h0; // @[Edges.scala 230:25]
  wire [127:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42]
  wire [127:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_75; // @[Monitor.scala 747:93]
  wire [127:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[127:1]}; // @[Monitor.scala 747:146]
  wire  _T_774 = io_in_d_valid & d_first_2 & _T_486; // @[Monitor.scala 779:71]
  wire [15:0] d_clr_1 = _d_first_T & d_first_2 & _T_486 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [142:0] _GEN_69 = _d_first_T & d_first_2 & _T_486 ? _d_sizes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 Monitor.scala 786:21]
  wire [15:0] _T_782 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0];
  wire  _T_792 = _GEN_83 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [15:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [15:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [127:0] d_sizes_clr_1 = _GEN_69[127:0];
  wire [127:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58]
  wire [127:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_812 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 10'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 10'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 10'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 10'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 16'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 64'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 128'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 10'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 10'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 10'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 10'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 16'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 128'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 10'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 10'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_98 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_98 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_T_98 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_106 & ~(_T_98 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_51 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_51 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_62 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_62 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_182 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(_T_330 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_284 & ~(_T_330 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(_T_364 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(_T_364 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_334 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(_T_364 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(_T_364 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_382 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(_T_64 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(_T_64 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(_T_228 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_430 & ~(_T_228 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_482 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_482 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_490 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_490 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_498 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_498 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_502 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_486 & ~(_T_502 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(_T_490 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(_T_490 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(_T_498 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_506 & ~(_T_498 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(_T_490 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(_T_490 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(_T_554 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_534 & ~(_T_554 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_563 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_563 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_563 & ~(_T_498 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_563 & ~(_T_498 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_580 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_580 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_580 & ~(_T_554 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_580 & ~(_T_554 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_598 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_598 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_598 & ~(_T_498 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_598 & ~(_T_498 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628 & ~(_T_629 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628 & ~(_T_629 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628 & ~(_T_637 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628 & ~(_T_637 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628 & ~(_T_641 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628 & ~(_T_641 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628 & ~(_T_645 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628 & ~(_T_645 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & ~(_T_653 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & ~(_T_653 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & ~(_T_661 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & ~(_T_661 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & ~(_T_665 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & ~(_T_665 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & ~(_T_673 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & ~(_T_673 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_682 & ~(_T_686 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_682 & ~(_T_686 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & ~(_T_705 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & ~(_T_705 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & same_cycle_resp & ~(_T_711 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & same_cycle_resp & ~(_T_711 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & same_cycle_resp & ~(_T_715 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & same_cycle_resp & ~(_T_715 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & ~same_cycle_resp & ~(_T_723 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & ~same_cycle_resp & ~(_T_723 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_693 & ~same_cycle_resp & ~(_T_727 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_693 & ~same_cycle_resp & ~(_T_727 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_737 & ~(_T_739 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_737 & ~(_T_739 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_748 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_748 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_774 & ~(_T_782[0] | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_774 & ~(_T_782[0] | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_774 & ~(_T_792 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_774 & ~(_T_792 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_812 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_812 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  source = _RAND_3[3:0];
  _RAND_4 = {4{`RANDOM}};
  address = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  d_first_counter = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  opcode_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  size_1 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  source_1 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  denied = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  inflight = _RAND_10[15:0];
  _RAND_11 = {2{`RANDOM}};
  inflight_opcodes = _RAND_11[63:0];
  _RAND_12 = {4{`RANDOM}};
  inflight_sizes = _RAND_12[127:0];
  _RAND_13 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  watchdog = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  inflight_1 = _RAND_16[15:0];
  _RAND_17 = {4{`RANDOM}};
  inflight_sizes_1 = _RAND_17[127:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[9:0];
  _RAND_19 = {1{`RANDOM}};
  watchdog_1 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLError_1(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [3:0]   auto_in_a_bits_size,
  input  [3:0]   auto_in_a_bits_source,
  input  [127:0] auto_in_a_bits_address,
  input  [3:0]   auto_in_a_bits_mask,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [2:0]   auto_in_d_bits_opcode,
  output [3:0]   auto_in_d_bits_size,
  output [3:0]   auto_in_d_bits_source,
  output         auto_in_d_bits_denied,
  output         auto_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [127:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  reg  idle; // @[Error.scala 44:23]
  reg [9:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle_1 = beatsLeft == 10'h0; // @[Arbiter.scala 88:28]
  reg [9:0] a_last_counter; // @[Edges.scala 228:27]
  wire  a_last_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [26:0] _a_last_beats1_decode_T_1 = 27'hfff << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [11:0] _a_last_beats1_decode_T_3 = ~_a_last_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [9:0] a_last_beats1_decode = _a_last_beats1_decode_T_3[11:2]; // @[Edges.scala 219:59]
  wire [9:0] a_last_beats1 = a_last_beats1_opdata ? a_last_beats1_decode : 10'h0; // @[Edges.scala 220:14]
  wire  a_last = a_last_counter == 10'h1 | a_last_beats1 == 10'h0; // @[Edges.scala 231:37]
  wire  da_valid = auto_in_a_valid & a_last & idle; // @[Error.scala 51:35]
  wire [1:0] _readys_T = {da_valid,1'h0}; // @[Cat.scala 30:58]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[package.scala 244:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[Arbiter.scala 16:61]
  wire  readys_1 = _readys_T_7[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle_1 ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_in_d_ready & allowed_1; // @[Arbiter.scala 123:31]
  reg [9:0] counter; // @[Edges.scala 228:27]
  wire [2:0] _GEN_4 = 3'h2 == auto_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_5 = 3'h3 == auto_in_a_bits_opcode ? 3'h1 : _GEN_4; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_6 = 3'h4 == auto_in_a_bits_opcode ? 3'h1 : _GEN_5; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_7 = 3'h5 == auto_in_a_bits_opcode ? 3'h2 : _GEN_6; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_8 = 3'h6 == auto_in_a_bits_opcode ? 3'h4 : _GEN_7; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] da_bits_opcode = 3'h7 == auto_in_a_bits_opcode ? 3'h4 : _GEN_8; // @[Error.scala 53:21 Error.scala 53:21]
  wire  beats1_opdata = da_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [9:0] beats1 = beats1_opdata ? a_last_beats1_decode : 10'h0; // @[Edges.scala 220:14]
  wire  da_last = counter == 10'h1 | beats1 == 10'h0; // @[Edges.scala 231:37]
  wire  in_a_ready = out_1_ready & da_last & idle | ~a_last; // @[Error.scala 50:46]
  wire  _a_last_T = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37]
  wire [9:0] a_last_counter1 = a_last_counter - 10'h1; // @[Edges.scala 229:28]
  wire  a_last_first = a_last_counter == 10'h0; // @[Edges.scala 230:25]
  wire  _T = out_1_ready & da_valid; // @[Decoupled.scala 40:37]
  wire [9:0] counter1 = counter - 10'h1; // @[Edges.scala 229:28]
  wire  da_first = counter == 10'h0; // @[Edges.scala 230:25]
  wire  _GEN_12 = _T & da_bits_opcode == 3'h4 ? 1'h0 : idle; // @[Error.scala 70:52 Error.scala 70:59 Error.scala 44:23]
  wire  latch = idle_1 & auto_in_d_ready; // @[Arbiter.scala 89:24]
  wire  earlyWinner_1 = readys_1 & da_valid; // @[Arbiter.scala 97:79]
  wire  _T_22 = ~da_valid; // @[Arbiter.scala 107:15]
  wire  muxStateEarly_1 = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_2 = state_1 & da_valid; // @[Mux.scala 27:72]
  wire  sink_ACancel_earlyValid = idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 50:33]
  wire [9:0] _GEN_17 = {{9'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [9:0] _beatsLeft_T_4 = beatsLeft - _GEN_17; // @[Arbiter.scala 113:52]
  TLMonitor_4 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  assign auto_in_a_ready = out_1_ready & da_last & idle | ~a_last; // @[Error.scala 50:46]
  assign auto_in_d_valid = idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2; // @[Arbiter.scala 125:29]
  assign auto_in_d_bits_opcode = muxStateEarly_1 ? da_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_size = muxStateEarly_1 ? auto_in_a_bits_size : 4'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_source = muxStateEarly_1 ? auto_in_a_bits_source : 4'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_denied = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  assign auto_in_d_bits_corrupt = muxStateEarly_1 & beats1_opdata; // @[Mux.scala 27:72]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = out_1_ready & da_last & idle | ~a_last; // @[Error.scala 50:46]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = idle_1 ? da_valid : _sink_ACancel_earlyValid_T_2; // @[Arbiter.scala 125:29]
  assign monitor_io_in_d_bits_opcode = muxStateEarly_1 ? da_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_size = muxStateEarly_1 ? auto_in_a_bits_size : 4'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_source = muxStateEarly_1 ? auto_in_a_bits_source : 4'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_denied = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  assign monitor_io_in_d_bits_corrupt = muxStateEarly_1 & beats1_opdata; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    idle <= reset | _GEN_12; // @[Error.scala 44:23 Error.scala 44:23]
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 10'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin // @[Arbiter.scala 113:23]
      if (earlyWinner_1) begin // @[Arbiter.scala 111:73]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          beatsLeft <= a_last_beats1_decode;
        end else begin
          beatsLeft <= 10'h0;
        end
      end else begin
        beatsLeft <= 10'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_last_counter <= 10'h0; // @[Edges.scala 228:27]
    end else if (_a_last_T) begin // @[Edges.scala 234:17]
      if (a_last_first) begin // @[Edges.scala 235:21]
        if (a_last_beats1_opdata) begin // @[Edges.scala 220:14]
          a_last_counter <= a_last_beats1_decode;
        end else begin
          a_last_counter <= 10'h0;
        end
      end else begin
        a_last_counter <= a_last_counter1;
      end
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin // @[Arbiter.scala 117:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 10'h0; // @[Edges.scala 228:27]
    end else if (_T) begin // @[Edges.scala 234:17]
      if (da_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          counter <= a_last_beats1_decode;
        end else begin
          counter <= 10'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(idle | da_first | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Error.scala:49 assert (idle || da_first) // we only send Grant, never GrantData => simplified flow control below\n"
            ); // @[Error.scala 49:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(idle | da_first | reset)) begin
          $fatal; // @[Error.scala 49:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~da_valid | earlyWinner_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~da_valid | earlyWinner_1 | reset)) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_22 | da_valid | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_22 | da_valid | reset)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  idle = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  beatsLeft = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  a_last_counter = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  state_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  counter = _RAND_4[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBusBypass(
  input         clock,
  input         reset,
  input         auto_node_out_out_a_ready,
  output        auto_node_out_out_a_valid,
  output [2:0]  auto_node_out_out_a_bits_opcode,
  output [2:0]  auto_node_out_out_a_bits_size,
  output [3:0]  auto_node_out_out_a_bits_source,
  output [31:0] auto_node_out_out_a_bits_address,
  output [3:0]  auto_node_out_out_a_bits_mask,
  output [31:0] auto_node_out_out_a_bits_data,
  output        auto_node_out_out_d_ready,
  input         auto_node_out_out_d_valid,
  input  [2:0]  auto_node_out_out_d_bits_opcode,
  input  [1:0]  auto_node_out_out_d_bits_param,
  input  [2:0]  auto_node_out_out_d_bits_size,
  input  [3:0]  auto_node_out_out_d_bits_source,
  input  [4:0]  auto_node_out_out_d_bits_sink,
  input         auto_node_out_out_d_bits_denied,
  input  [31:0] auto_node_out_out_d_bits_data,
  input         auto_node_out_out_d_bits_corrupt,
  output        auto_node_in_in_a_ready,
  input         auto_node_in_in_a_valid,
  input  [2:0]  auto_node_in_in_a_bits_opcode,
  input  [2:0]  auto_node_in_in_a_bits_size,
  input  [3:0]  auto_node_in_in_a_bits_source,
  input  [31:0] auto_node_in_in_a_bits_address,
  input  [3:0]  auto_node_in_in_a_bits_mask,
  input  [31:0] auto_node_in_in_a_bits_data,
  input         auto_node_in_in_d_ready,
  output        auto_node_in_in_d_valid,
  output [2:0]  auto_node_in_in_d_bits_opcode,
  output [1:0]  auto_node_in_in_d_bits_param,
  output [2:0]  auto_node_in_in_d_bits_size,
  output [3:0]  auto_node_in_in_d_bits_source,
  output [4:0]  auto_node_in_in_d_bits_sink,
  output        auto_node_in_in_d_bits_denied,
  output [31:0] auto_node_in_in_d_bits_data,
  output        auto_node_in_in_d_bits_corrupt,
  input         io_bypass
);
  wire  bar_clock; // @[BusBypass.scala 17:33]
  wire  bar_reset; // @[BusBypass.scala 17:33]
  wire  bar_auto_in_a_ready; // @[BusBypass.scala 17:33]
  wire  bar_auto_in_a_valid; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_in_a_bits_opcode; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_in_a_bits_size; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_in_a_bits_source; // @[BusBypass.scala 17:33]
  wire [31:0] bar_auto_in_a_bits_address; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_in_a_bits_mask; // @[BusBypass.scala 17:33]
  wire [31:0] bar_auto_in_a_bits_data; // @[BusBypass.scala 17:33]
  wire  bar_auto_in_d_ready; // @[BusBypass.scala 17:33]
  wire  bar_auto_in_d_valid; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_in_d_bits_opcode; // @[BusBypass.scala 17:33]
  wire [1:0] bar_auto_in_d_bits_param; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_in_d_bits_size; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_in_d_bits_source; // @[BusBypass.scala 17:33]
  wire [4:0] bar_auto_in_d_bits_sink; // @[BusBypass.scala 17:33]
  wire  bar_auto_in_d_bits_denied; // @[BusBypass.scala 17:33]
  wire [31:0] bar_auto_in_d_bits_data; // @[BusBypass.scala 17:33]
  wire  bar_auto_in_d_bits_corrupt; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_1_a_ready; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_1_a_valid; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_out_1_a_bits_opcode; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_out_1_a_bits_size; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_out_1_a_bits_source; // @[BusBypass.scala 17:33]
  wire [31:0] bar_auto_out_1_a_bits_address; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_out_1_a_bits_mask; // @[BusBypass.scala 17:33]
  wire [31:0] bar_auto_out_1_a_bits_data; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_1_d_ready; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_1_d_valid; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_out_1_d_bits_opcode; // @[BusBypass.scala 17:33]
  wire [1:0] bar_auto_out_1_d_bits_param; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_out_1_d_bits_size; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_out_1_d_bits_source; // @[BusBypass.scala 17:33]
  wire [4:0] bar_auto_out_1_d_bits_sink; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_1_d_bits_denied; // @[BusBypass.scala 17:33]
  wire [31:0] bar_auto_out_1_d_bits_data; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_1_d_bits_corrupt; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_0_a_ready; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_0_a_valid; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_out_0_a_bits_opcode; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_out_0_a_bits_size; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_out_0_a_bits_source; // @[BusBypass.scala 17:33]
  wire [127:0] bar_auto_out_0_a_bits_address; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_out_0_a_bits_mask; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_0_d_ready; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_0_d_valid; // @[BusBypass.scala 17:33]
  wire [2:0] bar_auto_out_0_d_bits_opcode; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_out_0_d_bits_size; // @[BusBypass.scala 17:33]
  wire [3:0] bar_auto_out_0_d_bits_source; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_0_d_bits_denied; // @[BusBypass.scala 17:33]
  wire  bar_auto_out_0_d_bits_corrupt; // @[BusBypass.scala 17:33]
  wire  bar_io_bypass; // @[BusBypass.scala 17:33]
  wire  error_clock; // @[BusBypass.scala 27:40]
  wire  error_reset; // @[BusBypass.scala 27:40]
  wire  error_auto_in_a_ready; // @[BusBypass.scala 27:40]
  wire  error_auto_in_a_valid; // @[BusBypass.scala 27:40]
  wire [2:0] error_auto_in_a_bits_opcode; // @[BusBypass.scala 27:40]
  wire [3:0] error_auto_in_a_bits_size; // @[BusBypass.scala 27:40]
  wire [3:0] error_auto_in_a_bits_source; // @[BusBypass.scala 27:40]
  wire [127:0] error_auto_in_a_bits_address; // @[BusBypass.scala 27:40]
  wire [3:0] error_auto_in_a_bits_mask; // @[BusBypass.scala 27:40]
  wire  error_auto_in_d_ready; // @[BusBypass.scala 27:40]
  wire  error_auto_in_d_valid; // @[BusBypass.scala 27:40]
  wire [2:0] error_auto_in_d_bits_opcode; // @[BusBypass.scala 27:40]
  wire [3:0] error_auto_in_d_bits_size; // @[BusBypass.scala 27:40]
  wire [3:0] error_auto_in_d_bits_source; // @[BusBypass.scala 27:40]
  wire  error_auto_in_d_bits_denied; // @[BusBypass.scala 27:40]
  wire  error_auto_in_d_bits_corrupt; // @[BusBypass.scala 27:40]
  TLBusBypassBar bar ( // @[BusBypass.scala 17:33]
    .clock(bar_clock),
    .reset(bar_reset),
    .auto_in_a_ready(bar_auto_in_a_ready),
    .auto_in_a_valid(bar_auto_in_a_valid),
    .auto_in_a_bits_opcode(bar_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(bar_auto_in_a_bits_size),
    .auto_in_a_bits_source(bar_auto_in_a_bits_source),
    .auto_in_a_bits_address(bar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(bar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(bar_auto_in_a_bits_data),
    .auto_in_d_ready(bar_auto_in_d_ready),
    .auto_in_d_valid(bar_auto_in_d_valid),
    .auto_in_d_bits_opcode(bar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(bar_auto_in_d_bits_param),
    .auto_in_d_bits_size(bar_auto_in_d_bits_size),
    .auto_in_d_bits_source(bar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(bar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(bar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(bar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(bar_auto_in_d_bits_corrupt),
    .auto_out_1_a_ready(bar_auto_out_1_a_ready),
    .auto_out_1_a_valid(bar_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(bar_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_size(bar_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(bar_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(bar_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_mask(bar_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_data(bar_auto_out_1_a_bits_data),
    .auto_out_1_d_ready(bar_auto_out_1_d_ready),
    .auto_out_1_d_valid(bar_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(bar_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_param(bar_auto_out_1_d_bits_param),
    .auto_out_1_d_bits_size(bar_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(bar_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_sink(bar_auto_out_1_d_bits_sink),
    .auto_out_1_d_bits_denied(bar_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_data(bar_auto_out_1_d_bits_data),
    .auto_out_1_d_bits_corrupt(bar_auto_out_1_d_bits_corrupt),
    .auto_out_0_a_ready(bar_auto_out_0_a_ready),
    .auto_out_0_a_valid(bar_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(bar_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_size(bar_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(bar_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(bar_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_mask(bar_auto_out_0_a_bits_mask),
    .auto_out_0_d_ready(bar_auto_out_0_d_ready),
    .auto_out_0_d_valid(bar_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(bar_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_size(bar_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(bar_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_denied(bar_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_corrupt(bar_auto_out_0_d_bits_corrupt),
    .io_bypass(bar_io_bypass)
  );
  TLError_1 error ( // @[BusBypass.scala 27:40]
    .clock(error_clock),
    .reset(error_reset),
    .auto_in_a_ready(error_auto_in_a_ready),
    .auto_in_a_valid(error_auto_in_a_valid),
    .auto_in_a_bits_opcode(error_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(error_auto_in_a_bits_size),
    .auto_in_a_bits_source(error_auto_in_a_bits_source),
    .auto_in_a_bits_address(error_auto_in_a_bits_address),
    .auto_in_a_bits_mask(error_auto_in_a_bits_mask),
    .auto_in_d_ready(error_auto_in_d_ready),
    .auto_in_d_valid(error_auto_in_d_valid),
    .auto_in_d_bits_opcode(error_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(error_auto_in_d_bits_size),
    .auto_in_d_bits_source(error_auto_in_d_bits_source),
    .auto_in_d_bits_denied(error_auto_in_d_bits_denied),
    .auto_in_d_bits_corrupt(error_auto_in_d_bits_corrupt)
  );
  assign auto_node_out_out_a_valid = bar_auto_out_1_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_node_out_out_a_bits_opcode = bar_auto_out_1_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_node_out_out_a_bits_size = bar_auto_out_1_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_node_out_out_a_bits_source = bar_auto_out_1_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_node_out_out_a_bits_address = bar_auto_out_1_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_node_out_out_a_bits_mask = bar_auto_out_1_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_node_out_out_a_bits_data = bar_auto_out_1_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_node_out_out_d_ready = bar_auto_out_1_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_node_in_in_a_ready = bar_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_valid = bar_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_bits_opcode = bar_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_bits_param = bar_auto_in_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_bits_size = bar_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_bits_source = bar_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_bits_sink = bar_auto_in_d_bits_sink; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_bits_denied = bar_auto_in_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_bits_data = bar_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_node_in_in_d_bits_corrupt = bar_auto_in_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign bar_clock = clock;
  assign bar_reset = reset;
  assign bar_auto_in_a_valid = auto_node_in_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bar_auto_in_a_bits_opcode = auto_node_in_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bar_auto_in_a_bits_size = auto_node_in_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bar_auto_in_a_bits_source = auto_node_in_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bar_auto_in_a_bits_address = auto_node_in_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bar_auto_in_a_bits_mask = auto_node_in_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bar_auto_in_a_bits_data = auto_node_in_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bar_auto_in_d_ready = auto_node_in_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bar_auto_out_1_a_ready = auto_node_out_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_valid = auto_node_out_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_bits_opcode = auto_node_out_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_bits_param = auto_node_out_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_bits_size = auto_node_out_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_bits_source = auto_node_out_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_bits_sink = auto_node_out_out_d_bits_sink; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_bits_denied = auto_node_out_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_bits_data = auto_node_out_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_1_d_bits_corrupt = auto_node_out_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bar_auto_out_0_a_ready = error_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign bar_auto_out_0_d_valid = error_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign bar_auto_out_0_d_bits_opcode = error_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign bar_auto_out_0_d_bits_size = error_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign bar_auto_out_0_d_bits_source = error_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign bar_auto_out_0_d_bits_denied = error_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign bar_auto_out_0_d_bits_corrupt = error_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign bar_io_bypass = io_bypass; // @[BusBypass.scala 44:26]
  assign error_clock = clock;
  assign error_reset = reset;
  assign error_auto_in_a_valid = bar_auto_out_0_a_valid; // @[LazyModule.scala 298:16]
  assign error_auto_in_a_bits_opcode = bar_auto_out_0_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign error_auto_in_a_bits_size = bar_auto_out_0_a_bits_size; // @[LazyModule.scala 298:16]
  assign error_auto_in_a_bits_source = bar_auto_out_0_a_bits_source; // @[LazyModule.scala 298:16]
  assign error_auto_in_a_bits_address = bar_auto_out_0_a_bits_address; // @[LazyModule.scala 298:16]
  assign error_auto_in_a_bits_mask = bar_auto_out_0_a_bits_mask; // @[LazyModule.scala 298:16]
  assign error_auto_in_d_ready = bar_auto_out_0_d_ready; // @[LazyModule.scala 298:16]
endmodule
module TLMonitor_5(
  input        clock,
  input        reset,
  input        io_in_d_valid,
  input  [2:0] io_in_d_bits_opcode,
  input  [1:0] io_in_d_bits_param,
  input  [2:0] io_in_d_bits_size,
  input        io_in_d_bits_source,
  input        io_in_d_bits_denied,
  input        io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _T_677 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9]
  wire  _T_681 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_685 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_689 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_693 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_697 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_701 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_712 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_716 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_729 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_749 = _T_697 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_758 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_775 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_793 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg  source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_1648 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_1649 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_1653 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_1657 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_1661 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_1669 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [3:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [2:0] _GEN_86 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_86}; // @[Monitor.scala 634:69]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [15:0] _GEN_87 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_87 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152]
  wire [3:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [15:0] _GEN_90 = {{12'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91]
  wire [15:0] _a_size_lookup_T_6 = _GEN_90 & _a_opcode_lookup_T_5; // @[Monitor.scala 638:91]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144]
  wire  _T_1737 = io_in_d_valid & d_first_1 & ~_T_681; // @[Monitor.scala 671:71]
  wire [30:0] _GEN_93 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_93 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [30:0] _GEN_35 = _T_1737 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _T_1747 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_1766 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_1767 = io_in_d_bits_opcode == _GEN_60 | _T_1766; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_96 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_1771 = _GEN_96 == a_size_lookup; // @[Monitor.scala 691:36]
  wire [3:0] d_opcodes_clr = _GEN_35[3:0];
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [3:0] _inflight_opcodes_T_2 = inflight_opcodes & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [3:0] _inflight_sizes_T_2 = inflight_sizes & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [3:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [3:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [15:0] _GEN_101 = {{12'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93]
  wire [15:0] _c_size_lookup_T_6 = _GEN_101 & _a_opcode_lookup_T_5; // @[Monitor.scala 747:93]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146]
  wire  _T_1825 = io_in_d_valid & d_first_2 & _T_681; // @[Monitor.scala 779:71]
  wire [30:0] _GEN_80 = _T_1825 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_1843 = _GEN_96 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [3:0] d_opcodes_clr_1 = _GEN_80[3:0];
  wire [3:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [3:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [3:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_3 = d_first_counter_3 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 4'h0; // @[Edges.scala 230:25]
  wire  _T_1880 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_1881 = io_in_d_valid & d_first_3 & _T_1880; // @[Monitor.scala 829:38]
  wire  _T_1884 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = io_in_d_valid & d_first_3 & _T_1880 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  d_set = _GEN_84[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (io_in_d_valid) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (io_in_d_valid & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (io_in_d_valid & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (io_in_d_valid & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (io_in_d_valid & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (io_in_d_valid & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 4'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (io_in_d_valid) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 4'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (io_in_d_valid) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= inflight_2 | d_set; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 4'h0; // @[Edges.scala 228:27]
    end else if (io_in_d_valid) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 4'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_677 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_677 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_source_ok_T_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_source_ok_T_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_T_685 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_T_685 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_T_689 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_T_689 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_T_693 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_T_693 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_T_697 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_681 & ~(_T_697 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_source_ok_T_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_source_ok_T_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_T_685 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_T_685 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_T_712 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_T_712 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_T_716 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_T_716 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_T_693 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_701 & ~(_T_693 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_source_ok_T_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_source_ok_T_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_T_685 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_T_685 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_T_712 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_T_712 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_T_716 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_T_716 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_T_749 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_729 & ~(_T_749 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_758 & ~(_source_ok_T_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_758 & ~(_source_ok_T_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_758 & ~(_T_689 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_758 & ~(_T_689 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_758 & ~(_T_693 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_758 & ~(_T_693 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_775 & ~(_source_ok_T_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_775 & ~(_source_ok_T_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_775 & ~(_T_689 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_775 & ~(_T_689 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_775 & ~(_T_749 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_775 & ~(_T_749 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_793 & ~(_source_ok_T_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_793 & ~(_source_ok_T_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_793 & ~(_T_689 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_793 & ~(_T_689 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_793 & ~(_T_693 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_793 & ~(_T_693 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1648 & ~(_T_1649 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1648 & ~(_T_1649 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1648 & ~(_T_1653 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1648 & ~(_T_1653 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1648 & ~(_T_1657 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1648 & ~(_T_1657 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1648 & ~(_T_1661 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1648 & ~(_T_1661 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1648 & ~(_T_1669 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1648 & ~(_T_1669 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1737 & ~(_T_1747 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1737 & ~(_T_1747 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1737 & ~(_T_1767 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1737 & ~(_T_1767 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1737 & ~(_T_1771 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1737 & ~(_T_1771 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1825 & ~(_T_1747 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1825 & ~(_T_1747 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1825 & ~(_T_1843 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1825 & ~(_T_1843 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1881 & ~(_T_1884 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLink.scala:70:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1881 & ~(_T_1884 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  d_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param_1 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  size_1 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  denied = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  inflight_opcodes = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  inflight_sizes = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  inflight_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_12[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_6(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [5:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [3:0]  io_in_a_bits_mask,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [2:0]  io_in_c_bits_size,
  input  [5:0]  io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [5:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input         io_in_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [255:0] _RAND_19;
  reg [255:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [255:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_86 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire [31:0] _T_180 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_181 = {1'b0,$signed(_T_180)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_183 = $signed(_T_181) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_184 = $signed(_T_183) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_185 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_186 = {1'b0,$signed(_T_185)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_188 = $signed(_T_186) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_189 = $signed(_T_188) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_190 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_191 = {1'b0,$signed(_T_190)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_193 = $signed(_T_191) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_194 = $signed(_T_193) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_195 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_196 = {1'b0,$signed(_T_195)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_198 = $signed(_T_196) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_199 = $signed(_T_198) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_200 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_201 = {1'b0,$signed(_T_200)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_203 = $signed(_T_201) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_204 = $signed(_T_203) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_211 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_214 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_215 = {1'b0,$signed(_T_214)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_217 = $signed(_T_215) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_218 = $signed(_T_217) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_219 = _T_211 & _T_218; // @[Parameters.scala 670:56]
  wire  _T_222 = source_ok & _T_219; // @[Monitor.scala 82:72]
  wire  _T_277 = _source_ok_T_1 & _T_211; // @[Mux.scala 27:72]
  wire  _T_330 = _T_218 | _T_184 | _T_189 | _T_194 | _T_199 | _T_204; // @[Parameters.scala 671:42]
  wire  _T_333 = _T_277 & _T_330; // @[Monitor.scala 83:78]
  wire  _T_347 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [3:0] _T_351 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_352 = _T_351 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_360 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_593 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_606 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_709 = _T_211 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_720 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_724 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_732 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_834 = source_ok & _T_709; // @[Monitor.scala 115:71]
  wire  _T_852 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_968 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_969 = io_in_a_bits_mask & _T_968; // @[Monitor.scala 127:31]
  wire  _T_970 = _T_969 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_974 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_1036 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_1074 = _T_1036 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_1076 = source_ok & _T_1074; // @[Monitor.scala 131:74]
  wire  _T_1086 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_1094 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_1206 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_1214 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1326 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1338 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1342 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1346 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_1350 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_1354 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1358 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1362 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1373 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_1377 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_1390 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1410 = _T_1358 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1419 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1436 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1454 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _source_ok_T_109 = io_in_c_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_115 = io_in_c_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_121 = io_in_c_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_127 = io_in_c_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_133 = io_in_c_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_139 = io_in_c_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_145 = io_in_c_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_151 = io_in_c_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_2 = _source_ok_T_109 | _source_ok_T_115 | _source_ok_T_121 | _source_ok_T_127 | _source_ok_T_133 |
    _source_ok_T_139 | _source_ok_T_145 | _source_ok_T_151; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_7 = 13'h3f << io_in_c_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask_2 = ~_is_aligned_mask_T_7[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_87 = {{26'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T_2 = io_in_c_bits_address & _GEN_87; // @[Edges.scala 20:16]
  wire  is_aligned_2 = _is_aligned_T_2 == 32'h0; // @[Edges.scala 20:24]
  wire [31:0] _address_ok_T_34 = io_in_c_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_35 = {1'b0,$signed(_address_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_37 = $signed(_address_ok_T_35) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_38 = $signed(_address_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_39 = io_in_c_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_40 = {1'b0,$signed(_address_ok_T_39)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_42 = $signed(_address_ok_T_40) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_43 = $signed(_address_ok_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_44 = io_in_c_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_45 = {1'b0,$signed(_address_ok_T_44)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_47 = $signed(_address_ok_T_45) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_48 = $signed(_address_ok_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_49 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_50 = {1'b0,$signed(_address_ok_T_49)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_52 = $signed(_address_ok_T_50) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_53 = $signed(_address_ok_T_52) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_54 = io_in_c_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_55 = {1'b0,$signed(_address_ok_T_54)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_57 = $signed(_address_ok_T_55) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_58 = $signed(_address_ok_T_57) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _address_ok_T_62 = _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 | _address_ok_T_58; // @[Parameters.scala 598:92]
  wire [31:0] _address_ok_T_63 = io_in_c_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_64 = {1'b0,$signed(_address_ok_T_63)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_66 = $signed(_address_ok_T_64) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_67 = $signed(_address_ok_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  wire  address_ok_1 = _address_ok_T_62 | _address_ok_T_67; // @[Parameters.scala 622:64]
  wire  _T_2224 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  wire  _T_2231 = io_in_c_bits_size >= 3'h2; // @[Monitor.scala 245:30]
  wire  _T_2238 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  wire  _T_2246 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  wire  _T_2264 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  wire  _T_2357 = io_in_c_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_2365 = _T_2357 & _address_ok_T_67; // @[Parameters.scala 670:56]
  wire  _T_2368 = source_ok_2 & _T_2365; // @[Monitor.scala 260:78]
  wire  _T_2423 = _source_ok_T_109 & _T_2357; // @[Mux.scala 27:72]
  wire  _T_2476 = _address_ok_T_67 | _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 |
    _address_ok_T_58; // @[Parameters.scala 671:42]
  wire  _T_2479 = _T_2423 & _T_2476; // @[Monitor.scala 261:78]
  wire  _T_2501 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  wire  _T_2734 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  wire  _T_2744 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  wire  _T_2752 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  wire  _T_2766 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  wire  sink_ok_1 = io_in_e_bits_sink < 1'h1; // @[Monitor.scala 364:31]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [5:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_2788 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_2789 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_2793 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_2797 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_2801 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_2805 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [5:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_2812 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_2813 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_2817 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_2821 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_2825 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_2833 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  wire  _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  wire [3:0] c_first_beats1_decode = is_aligned_mask_2[5:2]; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  reg [3:0] c_first_counter; // @[Edges.scala 228:27]
  wire [3:0] c_first_counter1 = c_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  c_first = c_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [2:0] size_3; // @[Monitor.scala 514:22]
  reg [5:0] source_3; // @[Monitor.scala 515:22]
  reg [31:0] address_2; // @[Monitor.scala 516:22]
  wire  _T_2864 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  wire  _T_2865 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  wire  _T_2869 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  wire  _T_2873 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  wire  _T_2877 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  wire  _T_2881 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  reg [63:0] inflight; // @[Monitor.scala 611:27]
  reg [255:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [255:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [7:0] _GEN_88 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [8:0] _a_opcode_lookup_T = {{1'd0}, _GEN_88}; // @[Monitor.scala 634:69]
  wire [255:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [255:0] _GEN_89 = {{240'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [255:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_89; // @[Monitor.scala 634:97]
  wire [255:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[255:1]}; // @[Monitor.scala 634:152]
  wire [255:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [255:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 638:91]
  wire [255:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[255:1]}; // @[Monitor.scala 638:144]
  wire  _T_2887 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [63:0] _a_set_wo_ready_T = 64'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 64'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_2890 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [7:0] _GEN_94 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [8:0] _a_opcodes_set_T = {{1'd0}, _GEN_94}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [514:0] _GEN_95 = {{511'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [514:0] _a_opcodes_set_T_1 = _GEN_95 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [514:0] _GEN_97 = {{511'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [514:0] _a_sizes_set_T_1 = _GEN_97 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [63:0] _T_2892 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_2894 = ~_T_2892[0]; // @[Monitor.scala 658:17]
  wire [63:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 64'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [514:0] _GEN_31 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 515'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [514:0] _GEN_32 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 515'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_2898 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_2900 = ~_T_1342; // @[Monitor.scala 671:74]
  wire  _T_2901 = io_in_d_valid & d_first_1 & ~_T_1342; // @[Monitor.scala 671:71]
  wire [63:0] _d_clr_wo_ready_T = 64'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [526:0] _GEN_99 = {{511'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [526:0] _d_opcodes_clr_T_5 = _GEN_99 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [63:0] d_clr = _d_first_T & d_first_1 & _T_2900 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [526:0] _GEN_35 = _d_first_T & d_first_1 & _T_2900 ? _d_opcodes_clr_T_5 : 527'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_2887 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [63:0] _T_2911 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_2913 = _T_2911[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_2918 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_2919 = io_in_d_bits_opcode == _GEN_44 | _T_2918; // @[Monitor.scala 685:77]
  wire  _T_2923 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_2930 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_2931 = io_in_d_bits_opcode == _GEN_60 | _T_2930; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_102 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_2935 = _GEN_102 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_2945 = _T_2898 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_2900; // @[Monitor.scala 694:116]
  wire  _T_2946 = ~io_in_d_ready; // @[Monitor.scala 695:15]
  wire  _T_2947 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_2954 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [63:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [63:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [63:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [255:0] a_opcodes_set = _GEN_31[255:0];
  wire [255:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [255:0] d_opcodes_clr = _GEN_35[255:0];
  wire [255:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [255:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [255:0] a_sizes_set = _GEN_32[255:0];
  wire [255:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [255:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_2963 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [63:0] inflight_1; // @[Monitor.scala 723:35]
  reg [255:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] c_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] c_first_counter1_1 = c_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  c_first_1 = c_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [255:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [255:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 747:93]
  wire [255:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[255:1]}; // @[Monitor.scala 747:146]
  wire  _T_2973 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  _T_2974 = io_in_c_valid & c_first_1 & _T_2973; // @[Monitor.scala 756:37]
  wire [63:0] _c_set_wo_ready_T = 64'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] c_set_wo_ready = io_in_c_valid & c_first_1 & _T_2973 ? _c_set_wo_ready_T : 64'h0; // @[Monitor.scala 756:71 Monitor.scala 757:22]
  wire  _T_2980 = _c_first_T & c_first_1 & _T_2973; // @[Monitor.scala 760:38]
  wire [3:0] _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  wire [3:0] _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 4'h1; // @[Monitor.scala 763:59]
  wire [7:0] _GEN_109 = {io_in_c_bits_source, 2'h0}; // @[Monitor.scala 764:79]
  wire [8:0] _c_opcodes_set_T = {{1'd0}, _GEN_109}; // @[Monitor.scala 764:79]
  wire [3:0] c_sizes_set_interm = _c_first_T & c_first_1 & _T_2973 ? _c_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 760:72 Monitor.scala 763:28]
  wire [514:0] _GEN_112 = {{511'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  wire [514:0] _c_sizes_set_T_1 = _GEN_112 << _c_opcodes_set_T; // @[Monitor.scala 765:52]
  wire [63:0] _T_2981 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  wire  _T_2983 = ~_T_2981[0]; // @[Monitor.scala 766:17]
  wire [63:0] c_set = _c_first_T & c_first_1 & _T_2973 ? _c_set_wo_ready_T : 64'h0; // @[Monitor.scala 760:72 Monitor.scala 761:28]
  wire [514:0] _GEN_77 = _c_first_T & c_first_1 & _T_2973 ? _c_sizes_set_T_1 : 515'h0; // @[Monitor.scala 760:72 Monitor.scala 765:28]
  wire  _T_2987 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  wire  _T_2989 = io_in_d_valid & d_first_2 & _T_1342; // @[Monitor.scala 779:71]
  wire [63:0] d_clr_wo_ready_1 = io_in_d_valid & d_first_2 & _T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 779:89 Monitor.scala 780:22]
  wire [63:0] d_clr_1 = _d_first_T & d_first_2 & _T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [526:0] _GEN_80 = _d_first_T & d_first_2 & _T_1342 ? _d_opcodes_clr_T_5 : 527'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire  _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1 = _T_2974 & io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:88]
  wire [63:0] _T_2997 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire  _T_2999 = _T_2997[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  wire  _T_3003 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_3007 = _GEN_102 == c_size_lookup; // @[Monitor.scala 795:36]
  wire  _T_3016 = _T_2987 & c_first_1 & io_in_c_valid & _same_cycle_resp_T_8 & _T_1342; // @[Monitor.scala 799:116]
  wire  _T_3018 = _T_2946 | io_in_c_ready; // @[Monitor.scala 800:32]
  wire  _T_3022 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  wire  _T_3023 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  wire [63:0] _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  wire [63:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [63:0] _inflight_T_5 = _inflight_T_3 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [255:0] d_opcodes_clr_1 = _GEN_80[255:0];
  wire [255:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [255:0] c_sizes_set = _GEN_77[255:0];
  wire [255:0] _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  wire [255:0] _inflight_sizes_T_5 = _inflight_sizes_T_3 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_3032 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [3:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_3 = d_first_counter_3 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 4'h0; // @[Edges.scala 230:25]
  wire  _T_3044 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_3045 = _d_first_T & d_first_3 & _T_3044; // @[Monitor.scala 829:38]
  wire  _T_3048 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = _d_first_T & d_first_3 & _T_3044 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  _T_3052 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _e_clr_T = 2'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  wire  d_set = _GEN_84[0];
  wire  _T_3056 = (d_set | inflight_2) >> io_in_e_bits_sink; // @[Monitor.scala 837:35]
  wire [1:0] _GEN_85 = _T_3052 ? _e_clr_T : 2'h0; // @[Monitor.scala 835:73 Monitor.scala 836:13]
  wire  e_clr = _GEN_85[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 4'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      opcode_3 <= io_in_c_bits_opcode; // @[Monitor.scala 525:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      param_3 <= io_in_c_bits_param; // @[Monitor.scala 526:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      size_3 <= io_in_c_bits_size; // @[Monitor.scala 527:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      source_3 <= io_in_c_bits_source; // @[Monitor.scala 528:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      address_2 <= io_in_c_bits_address; // @[Monitor.scala 529:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 64'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 256'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 256'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 64'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 256'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first_1) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 4'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_c_first_T | _d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= (inflight_2 | d_set) & ~e_clr; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 4'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1326 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1326 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1338 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1338 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1358 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1358 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1373 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1373 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1377 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1377 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1373 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1373 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1377 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1377 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1410 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1410 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2368 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2368 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2479 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2479 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid report param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2368 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2368 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2479 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2479 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid param (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channels carries invalid sink ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2789 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2789 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2793 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2793 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2797 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2797 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2801 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2805 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2813 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2813 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2817 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2817 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2821 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2821 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2825 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2825 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2833 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2833 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2865 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2865 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2869 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel param changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2869 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2873 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel size changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2873 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2877 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel source changed within multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2877 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2881 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel address changed with multibeat operation (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2881 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2890 & ~(_T_2894 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2890 & ~(_T_2894 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~(_T_2913 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~(_T_2913 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2919 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2919 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2923 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2923 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2931 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2931 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2935 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2935 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2945 & ~(_T_2947 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2945 & ~(_T_2947 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2954 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2954 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2963 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2963 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2980 & ~(_T_2983 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel re-used a source ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2980 & ~(_T_2983 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & ~(_T_2999 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & ~(_T_2999 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & same_cycle_resp_1 & ~(_T_3003 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & same_cycle_resp_1 & ~(_T_3003 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & ~same_cycle_resp_1 & ~(_T_3007 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & ~same_cycle_resp_1 & ~(_T_3007 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3016 & ~(_T_3018 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3016 & ~(_T_3018 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3022 & ~(_T_3023 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3022 & ~(_T_3023 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_3032 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_3032 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3045 & ~(_T_3048 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLink.scala:71:16)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3045 & ~(_T_3048 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3052 & ~(_T_3056 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChipLink.scala:71:16)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3052 & ~(_T_3056 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  c_first_counter = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  opcode_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  param_3 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  size_3 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  source_3 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  address_2 = _RAND_17[31:0];
  _RAND_18 = {2{`RANDOM}};
  inflight = _RAND_18[63:0];
  _RAND_19 = {8{`RANDOM}};
  inflight_opcodes = _RAND_19[255:0];
  _RAND_20 = {8{`RANDOM}};
  inflight_sizes = _RAND_20[255:0];
  _RAND_21 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  watchdog = _RAND_23[31:0];
  _RAND_24 = {2{`RANDOM}};
  inflight_1 = _RAND_24[63:0];
  _RAND_25 = {8{`RANDOM}};
  inflight_sizes_1 = _RAND_25[255:0];
  _RAND_26 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  watchdog_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inflight_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_30[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StuckSnooper(
  input         clock,
  input         reset,
  output        auto_in_1_a_ready,
  input         auto_in_1_a_valid,
  input  [2:0]  auto_in_1_a_bits_opcode,
  input  [2:0]  auto_in_1_a_bits_param,
  input  [2:0]  auto_in_1_a_bits_size,
  input  [5:0]  auto_in_1_a_bits_source,
  input  [31:0] auto_in_1_a_bits_address,
  input  [3:0]  auto_in_1_a_bits_mask,
  input  [31:0] auto_in_1_a_bits_data,
  output        auto_in_1_c_ready,
  input         auto_in_1_c_valid,
  input  [2:0]  auto_in_1_c_bits_opcode,
  input  [2:0]  auto_in_1_c_bits_param,
  input  [2:0]  auto_in_1_c_bits_size,
  input  [5:0]  auto_in_1_c_bits_source,
  input  [31:0] auto_in_1_c_bits_address,
  input         auto_in_1_d_ready,
  output        auto_in_1_d_valid,
  output [2:0]  auto_in_1_d_bits_opcode,
  output [1:0]  auto_in_1_d_bits_param,
  output [2:0]  auto_in_1_d_bits_size,
  output [5:0]  auto_in_1_d_bits_source,
  output        auto_in_1_d_bits_denied,
  output [31:0] auto_in_1_d_bits_data,
  output        auto_in_1_e_ready,
  input         auto_in_1_e_valid,
  input         auto_in_1_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [2:0]  auto_out_a_bits_size,
  output [5:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [3:0]  auto_out_a_bits_mask,
  output [31:0] auto_out_a_bits_data,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [2:0]  auto_out_c_bits_size,
  output [5:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [2:0]  auto_out_d_bits_size,
  input  [5:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [31:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output        auto_out_e_bits_sink,
  input         io_bypass
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_1_clock; // @[Nodes.scala 24:25]
  wire  monitor_1_reset; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_1_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_1_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_1_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_1_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_1_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_1_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_e_ready; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_e_valid; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_e_bits_sink; // @[Nodes.scala 24:25]
  reg  bypass; // @[StuckSnooper.scala 41:25]
  reg [7:0] flight; // @[Edges.scala 294:25]
  reg [3:0] stall_counter; // @[Edges.scala 228:27]
  wire  stall_first = stall_counter == 4'h0; // @[Edges.scala 230:25]
  wire  stall = bypass != io_bypass & stall_first; // @[StuckSnooper.scala 46:40]
  wire  _bundleOut_0_a_valid_T = ~stall; // @[StuckSnooper.scala 50:20]
  wire  _bundleOut_0_a_valid_T_1 = bypass ? 1'h0 : auto_in_1_a_valid; // @[StuckSnooper.scala 50:33]
  wire  out_a_valid = ~stall & _bundleOut_0_a_valid_T_1; // @[StuckSnooper.scala 50:27]
  wire  _T = auto_out_a_ready & out_a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] out_a_bits_size = bypass ? 3'h0 : auto_in_1_a_bits_size; // @[StuckSnooper.scala 52:22]
  wire [12:0] _beats1_decode_T_1 = 13'h3f << out_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] beats1_decode = _beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire [2:0] out_a_bits_opcode = bypass ? 3'h0 : auto_in_1_a_bits_opcode; // @[StuckSnooper.scala 52:22]
  wire  beats1_opdata = ~out_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] counter; // @[Edges.scala 228:27]
  wire [3:0] counter1 = counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = counter == 4'h0; // @[Edges.scala 230:25]
  reg  divertprobes; // @[StuckSnooper.scala 61:31]
  wire  bypass_c = bypass | divertprobes; // @[StuckSnooper.scala 64:24]
  wire  out_c_valid = bypass_c ? 1'h0 : auto_in_1_c_valid; // @[StuckSnooper.scala 75:25]
  wire  _T_2 = auto_out_c_ready & out_c_valid; // @[Decoupled.scala 40:37]
  wire [2:0] out_c_bits_size = bypass_c ? 3'h0 : auto_in_1_c_bits_size; // @[StuckSnooper.scala 77:24]
  wire [12:0] _beats1_decode_T_9 = 13'h3f << out_c_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_11 = ~_beats1_decode_T_9[5:0]; // @[package.scala 234:46]
  wire [3:0] beats1_decode_2 = _beats1_decode_T_11[5:2]; // @[Edges.scala 219:59]
  wire [2:0] out_c_bits_opcode = bypass_c ? 3'h4 : auto_in_1_c_bits_opcode; // @[StuckSnooper.scala 77:24]
  wire  beats1_opdata_2 = out_c_bits_opcode[0]; // @[Edges.scala 101:36]
  wire [3:0] beats1_2 = beats1_opdata_2 ? beats1_decode_2 : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] counter_2; // @[Edges.scala 228:27]
  wire [3:0] counter1_2 = counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  c_first = counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire  c_last = counter_2 == 4'h1 | beats1_2 == 4'h0; // @[Edges.scala 231:37]
  wire  out_d_ready = bypass | auto_in_1_d_ready; // @[StuckSnooper.scala 54:23]
  wire  _T_3 = out_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _beats1_decode_T_13 = 13'h3f << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_15 = ~_beats1_decode_T_13[5:0]; // @[package.scala 234:46]
  wire [3:0] beats1_decode_3 = _beats1_decode_T_15[5:2]; // @[Edges.scala 219:59]
  wire  beats1_opdata_3 = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [3:0] beats1_3 = beats1_opdata_3 ? beats1_decode_3 : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] counter_3; // @[Edges.scala 228:27]
  wire [3:0] counter1_3 = counter_3 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = counter_3 == 4'h0; // @[Edges.scala 230:25]
  wire  d_last = counter_3 == 4'h1 | beats1_3 == 4'h0; // @[Edges.scala 231:37]
  wire  out_e_valid = bypass_c ? 1'h0 : auto_in_1_e_valid; // @[StuckSnooper.scala 81:25]
  wire  done_4 = auto_out_e_ready & out_e_valid; // @[Decoupled.scala 40:37]
  wire  c_request = out_c_bits_opcode[2] & out_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  c_response = ~out_c_bits_opcode[2] | ~out_c_bits_opcode[1]; // @[Edges.scala 81:41]
  wire  d_request = auto_out_d_bits_opcode[2] & ~auto_out_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  inc_hi_hi_hi = _T & a_first; // @[Edges.scala 309:28]
  wire  inc_lo_hi = _T_2 & c_first & c_request; // @[Edges.scala 311:39]
  wire  inc_hi_hi_lo = _T_3 & d_first & d_request; // @[Edges.scala 312:39]
  wire [4:0] inc = {inc_hi_hi_hi,inc_hi_hi_lo,1'h0,inc_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire  dec_lo_hi = _T_2 & c_last & c_response; // @[Edges.scala 318:38]
  wire  dec_hi_hi_lo = _T_3 & d_last; // @[Edges.scala 319:28]
  wire [4:0] dec = {1'h0,dec_hi_hi_lo,1'h0,dec_lo_hi,done_4}; // @[Cat.scala 30:58]
  wire [1:0] _next_flight_T_5 = inc[0] + inc[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _next_flight_T_7 = inc[3] + inc[4]; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_7 = {{1'd0}, inc[2]}; // @[Bitwise.scala 47:55]
  wire [2:0] _next_flight_T_9 = _GEN_7 + _next_flight_T_7; // @[Bitwise.scala 47:55]
  wire [2:0] _next_flight_T_11 = _next_flight_T_5 + _next_flight_T_9[1:0]; // @[Bitwise.scala 47:55]
  wire [7:0] _GEN_8 = {{5'd0}, _next_flight_T_11}; // @[Edges.scala 323:30]
  wire [7:0] _next_flight_T_14 = flight + _GEN_8; // @[Edges.scala 323:30]
  wire [1:0] _next_flight_T_20 = dec[0] + dec[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _next_flight_T_22 = dec[3] + dec[4]; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_9 = {{1'd0}, dec[2]}; // @[Bitwise.scala 47:55]
  wire [2:0] _next_flight_T_24 = _GEN_9 + _next_flight_T_22; // @[Bitwise.scala 47:55]
  wire [2:0] _next_flight_T_26 = _next_flight_T_20 + _next_flight_T_24[1:0]; // @[Bitwise.scala 47:55]
  wire [7:0] _GEN_10 = {{5'd0}, _next_flight_T_26}; // @[Edges.scala 323:46]
  wire [7:0] next_flight = _next_flight_T_14 - _GEN_10; // @[Edges.scala 323:46]
  wire [3:0] stall_counter1 = stall_counter - 4'h1; // @[Edges.scala 229:28]
  wire  _bundleIn_0_a_ready_T_1 = _bundleOut_0_a_valid_T & auto_out_a_ready; // @[StuckSnooper.scala 48:27]
  wire  _bundleIn_1_a_ready_T_2 = ~bypass; // @[StuckSnooper.scala 49:45]
  wire  in1_a_ready = _bundleIn_0_a_ready_T_1 & ~bypass; // @[StuckSnooper.scala 49:42]
  wire  _divertprobes_T = in1_a_ready & auto_in_1_a_valid; // @[Decoupled.scala 40:37]
  wire  _bundleIn_1_bvalid_T = ~bypass_c; // @[StuckSnooper.scala 69:37]
  TLMonitor_5 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  TLMonitor_6 monitor_1 ( // @[Nodes.scala 24:25]
    .clock(monitor_1_clock),
    .reset(monitor_1_reset),
    .io_in_a_ready(monitor_1_io_in_a_ready),
    .io_in_a_valid(monitor_1_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_1_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_1_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_1_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_1_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_1_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_1_io_in_a_bits_mask),
    .io_in_c_ready(monitor_1_io_in_c_ready),
    .io_in_c_valid(monitor_1_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_1_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_1_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_1_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_1_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_1_io_in_c_bits_address),
    .io_in_d_ready(monitor_1_io_in_d_ready),
    .io_in_d_valid(monitor_1_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_1_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_1_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_1_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_1_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_1_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_1_io_in_d_bits_corrupt),
    .io_in_e_ready(monitor_1_io_in_e_ready),
    .io_in_e_valid(monitor_1_io_in_e_valid),
    .io_in_e_bits_sink(monitor_1_io_in_e_bits_sink)
  );
  assign auto_in_1_a_ready = _bundleIn_0_a_ready_T_1 & ~bypass; // @[StuckSnooper.scala 49:42]
  assign auto_in_1_c_ready = auto_out_c_ready & _bundleIn_1_bvalid_T; // @[StuckSnooper.scala 74:34]
  assign auto_in_1_d_valid = auto_out_d_valid & _bundleIn_1_a_ready_T_2; // @[StuckSnooper.scala 56:32]
  assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_e_ready = auto_out_e_ready & _bundleIn_1_bvalid_T; // @[StuckSnooper.scala 80:34]
  assign auto_out_a_valid = ~stall & _bundleOut_0_a_valid_T_1; // @[StuckSnooper.scala 50:27]
  assign auto_out_a_bits_opcode = bypass ? 3'h0 : auto_in_1_a_bits_opcode; // @[StuckSnooper.scala 52:22]
  assign auto_out_a_bits_param = bypass ? 3'h0 : auto_in_1_a_bits_param; // @[StuckSnooper.scala 52:22]
  assign auto_out_a_bits_size = bypass ? 3'h0 : auto_in_1_a_bits_size; // @[StuckSnooper.scala 52:22]
  assign auto_out_a_bits_source = bypass ? 6'h0 : auto_in_1_a_bits_source; // @[StuckSnooper.scala 52:22]
  assign auto_out_a_bits_address = bypass ? 32'h0 : auto_in_1_a_bits_address; // @[StuckSnooper.scala 52:22]
  assign auto_out_a_bits_mask = bypass ? 4'h0 : auto_in_1_a_bits_mask; // @[StuckSnooper.scala 52:22]
  assign auto_out_a_bits_data = bypass ? 32'h0 : auto_in_1_a_bits_data; // @[StuckSnooper.scala 52:22]
  assign auto_out_c_valid = bypass_c ? 1'h0 : auto_in_1_c_valid; // @[StuckSnooper.scala 75:25]
  assign auto_out_c_bits_opcode = bypass_c ? 3'h4 : auto_in_1_c_bits_opcode; // @[StuckSnooper.scala 77:24]
  assign auto_out_c_bits_param = bypass_c ? 3'h5 : auto_in_1_c_bits_param; // @[StuckSnooper.scala 77:24]
  assign auto_out_c_bits_size = bypass_c ? 3'h0 : auto_in_1_c_bits_size; // @[StuckSnooper.scala 77:24]
  assign auto_out_c_bits_source = bypass_c ? 6'h0 : auto_in_1_c_bits_source; // @[StuckSnooper.scala 77:24]
  assign auto_out_c_bits_address = bypass_c ? 32'h0 : auto_in_1_c_bits_address; // @[StuckSnooper.scala 77:24]
  assign auto_out_d_ready = bypass | auto_in_1_d_ready; // @[StuckSnooper.scala 54:23]
  assign auto_out_e_valid = bypass_c ? 1'h0 : auto_in_1_e_valid; // @[StuckSnooper.scala 81:25]
  assign auto_out_e_bits_sink = bypass_c ? 1'h0 : auto_in_1_e_bits_sink; // @[StuckSnooper.scala 83:24]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_d_valid = auto_out_d_valid & bypass; // @[StuckSnooper.scala 55:32]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source[0]; // @[Nodes.scala 1210:84 StuckSnooper.scala 57:16]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_a_ready = _bundleIn_0_a_ready_T_1 & ~bypass; // @[StuckSnooper.scala 49:42]
  assign monitor_1_io_in_a_valid = auto_in_1_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_a_bits_opcode = auto_in_1_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_a_bits_param = auto_in_1_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_a_bits_size = auto_in_1_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_a_bits_source = auto_in_1_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_a_bits_address = auto_in_1_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_a_bits_mask = auto_in_1_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_c_ready = auto_out_c_ready & _bundleIn_1_bvalid_T; // @[StuckSnooper.scala 74:34]
  assign monitor_1_io_in_c_valid = auto_in_1_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_c_bits_opcode = auto_in_1_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_c_bits_param = auto_in_1_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_c_bits_size = auto_in_1_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_c_bits_source = auto_in_1_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_c_bits_address = auto_in_1_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_d_ready = auto_in_1_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_d_valid = auto_out_d_valid & _bundleIn_1_a_ready_T_2; // @[StuckSnooper.scala 56:32]
  assign monitor_1_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_1_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_1_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_1_io_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_1_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_1_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_1_io_in_e_ready = auto_out_e_ready & _bundleIn_1_bvalid_T; // @[StuckSnooper.scala 80:34]
  assign monitor_1_io_in_e_valid = auto_in_1_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_1_io_in_e_bits_sink = auto_in_1_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  always @(posedge clock) begin
    if (reset) begin // @[StuckSnooper.scala 41:25]
      bypass <= io_bypass; // @[StuckSnooper.scala 41:25]
    end else if (next_flight == 8'h0) begin // @[StuckSnooper.scala 45:36]
      bypass <= io_bypass; // @[StuckSnooper.scala 45:45]
    end
    if (reset) begin // @[Edges.scala 294:25]
      flight <= 8'h0; // @[Edges.scala 294:25]
    end else begin
      flight <= next_flight; // @[Edges.scala 324:12]
    end
    if (reset) begin // @[Edges.scala 228:27]
      stall_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T) begin // @[Edges.scala 234:17]
      if (stall_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          stall_counter <= beats1_decode;
        end else begin
          stall_counter <= 4'h0;
        end
      end else begin
        stall_counter <= stall_counter1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          counter <= beats1_decode;
        end else begin
          counter <= 4'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    divertprobes <= reset | divertprobes & ~(_divertprobes_T & (auto_in_1_a_bits_opcode == 3'h6 |
      auto_in_1_a_bits_opcode == 3'h7)); // @[StuckSnooper.scala 61:31 StuckSnooper.scala 61:31 StuckSnooper.scala 62:18]
    if (reset) begin // @[Edges.scala 228:27]
      counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T_2) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata_2) begin // @[Edges.scala 220:14]
          counter_2 <= beats1_decode_2;
        end else begin
          counter_2 <= 4'h0;
        end
      end else begin
        counter_2 <= counter1_2;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter_3 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T_3) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata_3) begin // @[Edges.scala 220:14]
          counter_3 <= beats1_decode_3;
        end else begin
          counter_3 <= 4'h0;
        end
      end else begin
        counter_3 <= counter1_3;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bypass = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  flight = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  stall_counter = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  counter = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  divertprobes = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  counter_2 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  counter_3 = _RAND_6[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_7(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [3:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [3:0]  io_in_a_bits_mask,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [3:0]  io_in_d_bits_source,
  input  [4:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = ~io_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | io_in_a_bits_source[3]; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_34 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_60 = 3'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48]
  wire [31:0] _T_62 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_63 = {1'b0,$signed(_T_62)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_65 = $signed(_T_63) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_66 = $signed(_T_65) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_77 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_78 = {1'b0,$signed(_T_77)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_80 = $signed(_T_78) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_81 = $signed(_T_80) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_82 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_83 = {1'b0,$signed(_T_82)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_85 = $signed(_T_83) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_86 = $signed(_T_85) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_90 = _T_66 | _T_71 | _T_76 | _T_81 | _T_86; // @[Parameters.scala 671:42]
  wire  _T_91 = _T_60 & _T_90; // @[Parameters.scala 670:56]
  wire  _T_94 = source_ok & _T_91; // @[Monitor.scala 82:72]
  wire [32:0] _T_120 = $signed(_T_78) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _T_121 = $signed(_T_120) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_124 = _T_66 | _T_71 | _T_76 | _T_121; // @[Parameters.scala 671:42]
  wire [3:0] _T_145 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_146 = _T_145 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_154 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_278 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_301 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_327 = _T_301 & _T_124; // @[Parameters.scala 670:56]
  wire  _T_342 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_350 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_398 = source_ok & _T_327; // @[Monitor.scala 115:71]
  wire  _T_416 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_478 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_479 = io_in_a_bits_mask & _T_478; // @[Monitor.scala 127:31]
  wire  _T_480 = _T_479 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_484 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_504 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_530 = _T_504 & _T_124; // @[Parameters.scala 670:56]
  wire  _T_532 = source_ok & _T_530; // @[Monitor.scala 131:74]
  wire  _T_550 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_616 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_686 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_13 = ~io_in_d_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_13 | io_in_d_bits_source[3]; // @[Parameters.scala 1125:46]
  wire  _T_690 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_694 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_698 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_702 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_706 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_710 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_721 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_725 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_738 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_758 = _T_706 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_767 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_784 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_802 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [3:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_832 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_833 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_841 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_845 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_849 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [3:0] source_1; // @[Monitor.scala 538:22]
  reg [4:0] sink; // @[Monitor.scala 539:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_856 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_857 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_861 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_865 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_869 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_873 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29]
  wire  _T_877 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [15:0] inflight; // @[Monitor.scala 611:27]
  reg [63:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [63:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69]
  wire [63:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [63:0] _GEN_73 = {{48'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[63:1]}; // @[Monitor.scala 634:152]
  wire [63:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [63:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91]
  wire [63:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[63:1]}; // @[Monitor.scala 638:144]
  wire  _T_883 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [15:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_886 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [15:0] _T_888 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_890 = ~_T_888[0]; // @[Monitor.scala 658:17]
  wire [15:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [130:0] _GEN_19 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [130:0] _GEN_20 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_894 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_896 = ~_T_690; // @[Monitor.scala 671:74]
  wire  _T_897 = io_in_d_valid & d_first_1 & ~_T_690; // @[Monitor.scala 671:71]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [15:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_690 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [15:0] d_clr = _d_first_T & d_first_1 & _T_896 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [142:0] _GEN_23 = _d_first_T & d_first_1 & _T_896 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_883 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [15:0] _T_907 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_909 = _T_907[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_914 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39]
  wire  _T_915 = io_in_d_bits_opcode == _GEN_32 | _T_914; // @[Monitor.scala 685:77]
  wire  _T_919 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_926 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_927 = io_in_d_bits_opcode == _GEN_48 | _T_926; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_931 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_941 = _T_894 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_896; // @[Monitor.scala 694:116]
  wire  _T_943 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_950 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [15:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [15:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [15:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [63:0] a_opcodes_set = _GEN_19[63:0];
  wire [63:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [63:0] d_opcodes_clr = _GEN_23[63:0];
  wire [63:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [63:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [63:0] a_sizes_set = _GEN_20[63:0];
  wire [63:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [63:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_959 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [15:0] inflight_1; // @[Monitor.scala 723:35]
  reg [63:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [63:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [63:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93]
  wire [63:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[63:1]}; // @[Monitor.scala 747:146]
  wire  _T_985 = io_in_d_valid & d_first_2 & _T_690; // @[Monitor.scala 779:71]
  wire [15:0] d_clr_1 = _d_first_T & d_first_2 & _T_690 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [142:0] _GEN_68 = _d_first_T & d_first_2 & _T_690 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire [15:0] _T_993 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_1003 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [15:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [15:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [63:0] d_opcodes_clr_1 = _GEN_68[63:0];
  wire [63:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [63:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_1028 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 16'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 64'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 64'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 16'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 64'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_94 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_94 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_146 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_146 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_T_94 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_T_94 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_T_146 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_154 & ~(_T_146 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(_T_327 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(_T_327 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_278 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(_T_398 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(_T_398 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_350 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(_T_398 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(_T_398 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(_T_480 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_416 & ~(_T_480 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(_T_532 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(_T_532 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_484 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(_T_532 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(_T_532 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_550 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(_T_398 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(_T_398 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(_T_342 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_616 & ~(_T_342 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_686 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_686 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_694 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_694 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_698 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_698 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_702 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_702 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_706 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_690 & ~(_T_706 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_694 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_694 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_721 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_725 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_725 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_702 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_710 & ~(_T_702 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_694 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_694 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_721 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_721 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_725 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_725 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_758 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_738 & ~(_T_758 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(_T_698 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(_T_698 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(_T_702 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_767 & ~(_T_702 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(_T_698 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(_T_698 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(_T_758 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_784 & ~(_T_758 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(_T_698 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(_T_698 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(_T_702 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_802 & ~(_T_702 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & ~(_T_833 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & ~(_T_833 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & ~(_T_841 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & ~(_T_841 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & ~(_T_845 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & ~(_T_845 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & ~(_T_849 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & ~(_T_849 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_857 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_857 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_861 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_861 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_865 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_865 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_869 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_869 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_873 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_873 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_856 & ~(_T_877 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_856 & ~(_T_877 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_886 & ~(_T_890 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_886 & ~(_T_890 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & ~(_T_909 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & ~(_T_909 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & same_cycle_resp & ~(_T_915 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & same_cycle_resp & ~(_T_915 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & same_cycle_resp & ~(_T_919 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & same_cycle_resp & ~(_T_919 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & ~same_cycle_resp & ~(_T_927 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & ~same_cycle_resp & ~(_T_927 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_897 & ~same_cycle_resp & ~(_T_931 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_897 & ~same_cycle_resp & ~(_T_931 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_941 & ~(_T_943 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_941 & ~(_T_943 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_950 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 8 (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_950 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_959 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_959 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_985 & ~(_T_993[0] | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_985 & ~(_T_993[0] | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_985 & ~(_T_1003 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLink.scala:66:13)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_985 & ~(_T_1003 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1028 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLink.scala:66:13)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1028 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  source = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  address = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  d_first_counter = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  opcode_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  param_1 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  sink = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight = _RAND_12[15:0];
  _RAND_13 = {2{`RANDOM}};
  inflight_opcodes = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_sizes = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  watchdog = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  inflight_1 = _RAND_18[15:0];
  _RAND_19 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  watchdog_1 = _RAND_21[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PartialInjector(
  input         clock,
  input         reset,
  input         io_i_last,
  output        io_o_last,
  output        io_i_ready,
  input         io_i_valid,
  input  [2:0]  io_i_bits_opcode,
  input  [2:0]  io_i_bits_param,
  input  [2:0]  io_i_bits_size,
  input  [3:0]  io_i_bits_source,
  input  [31:0] io_i_bits_address,
  input  [3:0]  io_i_bits_mask,
  input  [31:0] io_i_bits_data,
  input         io_o_ready,
  output        io_o_valid,
  output [2:0]  io_o_bits_opcode,
  output [2:0]  io_o_bits_param,
  output [2:0]  io_o_bits_size,
  output [3:0]  io_o_bits_source,
  output [31:0] io_o_bits_address,
  output [31:0] io_o_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] state; // @[Partial.scala 76:22]
  reg [31:0] shift; // @[Partial.scala 77:22]
  wire  full = state[3]; // @[Partial.scala 78:20]
  wire  partial = io_i_bits_opcode == 3'h1; // @[Partial.scala 79:26]
  reg  last; // @[Partial.scala 81:21]
  wire [7:0] mixed_lo_lo_hi = io_i_bits_data[7:0]; // @[Partial.scala 85:46]
  wire [7:0] mixed_lo_hi_hi = io_i_bits_data[15:8]; // @[Partial.scala 85:46]
  wire [7:0] mixed_hi_lo_hi = io_i_bits_data[23:16]; // @[Partial.scala 85:46]
  wire [7:0] mixed_hi_hi_hi = io_i_bits_data[31:24]; // @[Partial.scala 85:46]
  wire  mixed_lo_lo_lo = io_i_bits_mask[0]; // @[Partial.scala 86:24]
  wire  mixed_lo_hi_lo = io_i_bits_mask[1]; // @[Partial.scala 86:24]
  wire  mixed_hi_lo_lo = io_i_bits_mask[2]; // @[Partial.scala 86:24]
  wire  mixed_hi_hi_lo = io_i_bits_mask[3]; // @[Partial.scala 86:24]
  wire [35:0] mixed = {mixed_hi_hi_hi,mixed_hi_hi_lo,mixed_hi_lo_hi,mixed_hi_lo_lo,mixed_lo_hi_hi,mixed_lo_hi_lo,
    mixed_lo_lo_hi,mixed_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [5:0] _wide_T = {state, 2'h0}; // @[Partial.scala 88:42]
  wire [98:0] _GEN_11 = {{63'd0}, mixed}; // @[Partial.scala 88:32]
  wire [98:0] _wide_T_1 = _GEN_11 << _wide_T; // @[Partial.scala 88:32]
  wire [98:0] _GEN_12 = {{67'd0}, shift}; // @[Partial.scala 88:23]
  wire [98:0] wide = _GEN_12 | _wide_T_1; // @[Partial.scala 88:23]
  wire  _T_1 = ~last; // @[Partial.scala 92:34]
  wire  _GEN_0 = (io_i_last | full) & ~last ? 1'h0 : io_o_ready; // @[Partial.scala 92:41 Partial.scala 93:18 Partial.scala 64:8]
  wire  _T_3 = io_o_ready & io_o_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _state_T_1 = state + 4'h1; // @[Partial.scala 99:22]
  wire [66:0] _GEN_2 = full | last ? 67'h0 : wide[98:32]; // @[Partial.scala 100:27 Partial.scala 102:15 Partial.scala 98:13]
  wire [66:0] _GEN_3 = _T_3 ? _GEN_2 : {{35'd0}, shift}; // @[Partial.scala 97:24 Partial.scala 77:22]
  wire [98:0] _GEN_6 = partial ? wide : {{67'd0}, io_i_bits_data}; // @[Partial.scala 84:18 Partial.scala 89:12 Partial.scala 64:8]
  wire [66:0] _GEN_8 = partial ? _GEN_3 : {{35'd0}, shift}; // @[Partial.scala 84:18 Partial.scala 77:22]
  assign io_o_last = partial ? last : io_i_last; // @[Partial.scala 82:19]
  assign io_i_ready = partial ? _GEN_0 : io_o_ready; // @[Partial.scala 84:18 Partial.scala 64:8]
  assign io_o_valid = io_i_valid; // @[Partial.scala 64:8]
  assign io_o_bits_opcode = io_i_bits_opcode; // @[Partial.scala 64:8]
  assign io_o_bits_param = io_i_bits_param; // @[Partial.scala 64:8]
  assign io_o_bits_size = io_i_bits_size; // @[Partial.scala 64:8]
  assign io_o_bits_source = io_i_bits_source; // @[Partial.scala 64:8]
  assign io_o_bits_address = io_i_bits_address; // @[Partial.scala 64:8]
  assign io_o_bits_data = _GEN_6[31:0];
  always @(posedge clock) begin
    if (reset) begin // @[Partial.scala 76:22]
      state <= 4'h0; // @[Partial.scala 76:22]
    end else if (partial) begin // @[Partial.scala 84:18]
      if (_T_3) begin // @[Partial.scala 97:24]
        if (full | last) begin // @[Partial.scala 100:27]
          state <= 4'h0; // @[Partial.scala 101:15]
        end else begin
          state <= _state_T_1; // @[Partial.scala 99:13]
        end
      end
    end
    if (reset) begin // @[Partial.scala 77:22]
      shift <= 32'h0; // @[Partial.scala 77:22]
    end else begin
      shift <= _GEN_8[31:0];
    end
    if (reset) begin // @[Partial.scala 81:21]
      last <= 1'h0; // @[Partial.scala 81:21]
    end else if (partial) begin // @[Partial.scala 84:18]
      if (_T_3) begin // @[Partial.scala 97:24]
        last <= io_i_last & _T_1; // @[Partial.scala 104:12]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  shift = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  last = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask,
  output [31:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_param [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] ram_source [0:0]; // @[Decoupled.scala 218:16]
  wire [3:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_address [0:0]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] ram_mask [0:0]; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_data [0:0]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_14 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 249:27 Decoupled.scala 249:36]
  wire  do_enq = empty ? _GEN_14 : _do_enq_T; // @[Decoupled.scala 246:18]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 246:18 Decoupled.scala 248:14]
  assign ram_opcode_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = 1'h0;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_param_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_param_MPORT_data = 3'h0;
  assign ram_param_MPORT_addr = 1'h0;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = 1'h0;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_address_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = 1'h0;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_mask_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = 1'h0;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 245:25 Decoupled.scala 245:40 Decoupled.scala 240:16]
  assign io_deq_bits_opcode = empty ? io_enq_bits_opcode : ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_param = empty ? 3'h0 : ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_source = empty ? io_enq_bits_source : ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_address = empty ? io_enq_bits_address : ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_mask = empty ? io_enq_bits_mask : ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      if (empty) begin // @[Decoupled.scala 246:18]
        if (io_deq_ready) begin // @[Decoupled.scala 249:27]
          maybe_full <= 1'h0; // @[Decoupled.scala 249:36]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinkA(
  input         clock,
  input         reset,
  output        io_a_ready,
  input         io_a_valid,
  input  [2:0]  io_a_bits_opcode,
  input  [2:0]  io_a_bits_size,
  input  [3:0]  io_a_bits_source,
  input  [31:0] io_a_bits_address,
  input  [3:0]  io_a_bits_mask,
  input  [31:0] io_a_bits_data,
  input         io_q_ready,
  output        io_q_valid,
  output [31:0] io_q_bits_data,
  output        io_q_bits_last,
  output [6:0]  io_q_bits_beats
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inject_clock; // @[SinkA.scala 21:22]
  wire  inject_reset; // @[SinkA.scala 21:22]
  wire  inject_io_i_last; // @[SinkA.scala 21:22]
  wire  inject_io_o_last; // @[SinkA.scala 21:22]
  wire  inject_io_i_ready; // @[SinkA.scala 21:22]
  wire  inject_io_i_valid; // @[SinkA.scala 21:22]
  wire [2:0] inject_io_i_bits_opcode; // @[SinkA.scala 21:22]
  wire [2:0] inject_io_i_bits_param; // @[SinkA.scala 21:22]
  wire [2:0] inject_io_i_bits_size; // @[SinkA.scala 21:22]
  wire [3:0] inject_io_i_bits_source; // @[SinkA.scala 21:22]
  wire [31:0] inject_io_i_bits_address; // @[SinkA.scala 21:22]
  wire [3:0] inject_io_i_bits_mask; // @[SinkA.scala 21:22]
  wire [31:0] inject_io_i_bits_data; // @[SinkA.scala 21:22]
  wire  inject_io_o_ready; // @[SinkA.scala 21:22]
  wire  inject_io_o_valid; // @[SinkA.scala 21:22]
  wire [2:0] inject_io_o_bits_opcode; // @[SinkA.scala 21:22]
  wire [2:0] inject_io_o_bits_param; // @[SinkA.scala 21:22]
  wire [2:0] inject_io_o_bits_size; // @[SinkA.scala 21:22]
  wire [3:0] inject_io_o_bits_source; // @[SinkA.scala 21:22]
  wire [31:0] inject_io_o_bits_address; // @[SinkA.scala 21:22]
  wire [31:0] inject_io_o_bits_data; // @[SinkA.scala 21:22]
  wire  inject_io_i_q_clock; // @[Decoupled.scala 296:21]
  wire  inject_io_i_q_reset; // @[Decoupled.scala 296:21]
  wire  inject_io_i_q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  inject_io_i_q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] inject_io_i_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] inject_io_i_q_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [3:0] inject_io_i_q_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire [31:0] inject_io_i_q_io_enq_bits_address; // @[Decoupled.scala 296:21]
  wire [3:0] inject_io_i_q_io_enq_bits_mask; // @[Decoupled.scala 296:21]
  wire [31:0] inject_io_i_q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  inject_io_i_q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  inject_io_i_q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] inject_io_i_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] inject_io_i_q_io_deq_bits_param; // @[Decoupled.scala 296:21]
  wire [2:0] inject_io_i_q_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [3:0] inject_io_i_q_io_deq_bits_source; // @[Decoupled.scala 296:21]
  wire [31:0] inject_io_i_q_io_deq_bits_address; // @[Decoupled.scala 296:21]
  wire [3:0] inject_io_i_q_io_deq_bits_mask; // @[Decoupled.scala 296:21]
  wire [31:0] inject_io_i_q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  _inject_io_i_last_T = inject_io_i_ready & inject_io_i_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _inject_io_i_last_beats1_decode_T_1 = 13'h3f << inject_io_i_bits_size; // @[package.scala 234:77]
  wire [5:0] _inject_io_i_last_beats1_decode_T_3 = ~_inject_io_i_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] inject_io_i_last_beats1_decode = _inject_io_i_last_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  inject_io_i_last_beats1_opdata = ~inject_io_i_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [3:0] inject_io_i_last_beats1 = inject_io_i_last_beats1_opdata ? inject_io_i_last_beats1_decode : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] inject_io_i_last_counter; // @[Edges.scala 228:27]
  wire [3:0] inject_io_i_last_counter1 = inject_io_i_last_counter - 4'h1; // @[Edges.scala 229:28]
  wire  inject_io_i_last_first = inject_io_i_last_counter == 4'h0; // @[Edges.scala 230:25]
  wire  a_hasData = ~inject_io_o_bits_opcode[2]; // @[Edges.scala 91:28]
  wire  a_partial = inject_io_o_bits_opcode == 3'h1; // @[SinkA.scala 27:33]
  reg [1:0] state; // @[SinkA.scala 30:22]
  wire  _T = io_q_ready & io_q_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T = a_hasData ? 2'h3 : 2'h0; // @[SinkA.scala 40:37]
  wire  _T_4 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T_2 = ~inject_io_o_last ? 2'h3 : 2'h0; // @[SinkA.scala 41:37]
  wire [1:0] _GEN_1 = _T_4 ? _state_T_2 : state; // @[Conditional.scala 39:67 SinkA.scala 41:31 SinkA.scala 30:22]
  wire [1:0] _GEN_2 = _T_3 ? _state_T : _GEN_1; // @[Conditional.scala 39:67 SinkA.scala 40:31]
  wire [2:0] _GEN_7 = 4'h1 == inject_io_o_bits_source ? 3'h1 : 3'h0; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_8 = 4'h2 == inject_io_o_bits_source ? 3'h2 : _GEN_7; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_9 = 4'h3 == inject_io_o_bits_source ? 3'h3 : _GEN_8; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_10 = 4'h4 == inject_io_o_bits_source ? 3'h4 : _GEN_9; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_11 = 4'h5 == inject_io_o_bits_source ? 3'h5 : _GEN_10; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_12 = 4'h6 == inject_io_o_bits_source ? 3'h6 : _GEN_11; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_13 = 4'h7 == inject_io_o_bits_source ? 3'h7 : _GEN_12; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_14 = 4'h8 == inject_io_o_bits_source ? 3'h0 : _GEN_13; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_15 = 4'h9 == inject_io_o_bits_source ? 3'h1 : _GEN_14; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_16 = 4'ha == inject_io_o_bits_source ? 3'h2 : _GEN_15; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_17 = 4'hb == inject_io_o_bits_source ? 3'h3 : _GEN_16; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_18 = 4'hc == inject_io_o_bits_source ? 3'h4 : _GEN_17; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_19 = 4'hd == inject_io_o_bits_source ? 3'h5 : _GEN_18; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_20 = 4'he == inject_io_o_bits_source ? 3'h6 : _GEN_19; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] _GEN_21 = 4'hf == inject_io_o_bits_source ? 3'h7 : _GEN_20; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [15:0] header_hi_hi_hi = {{13'd0}, _GEN_21}; // @[Parameters.scala 80:35]
  wire [1:0] _GEN_30 = 4'h8 == inject_io_o_bits_source ? 2'h2 : 2'h1; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [1:0] _GEN_31 = 4'h9 == inject_io_o_bits_source ? 2'h2 : _GEN_30; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [1:0] _GEN_32 = 4'ha == inject_io_o_bits_source ? 2'h2 : _GEN_31; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [1:0] _GEN_33 = 4'hb == inject_io_o_bits_source ? 2'h2 : _GEN_32; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [1:0] _GEN_34 = 4'hc == inject_io_o_bits_source ? 2'h2 : _GEN_33; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [1:0] _GEN_35 = 4'hd == inject_io_o_bits_source ? 2'h2 : _GEN_34; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [1:0] _GEN_36 = 4'he == inject_io_o_bits_source ? 2'h2 : _GEN_35; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [1:0] _GEN_37 = 4'hf == inject_io_o_bits_source ? 2'h2 : _GEN_36; // @[Parameters.scala 80:35 Parameters.scala 80:35]
  wire [2:0] header_hi_hi_lo = {{1'd0}, _GEN_37}; // @[Parameters.scala 80:35]
  wire [3:0] header_hi_lo = {{1'd0}, inject_io_o_bits_size}; // @[Parameters.scala 80:35]
  wire [2:0] header_lo_hi_hi = inject_io_o_bits_param; // @[Parameters.scala 80:35]
  wire [2:0] header_lo_hi_lo = inject_io_o_bits_opcode; // @[Parameters.scala 80:35]
  wire [31:0] header = {header_hi_hi_hi,header_hi_hi_lo,header_hi_lo,header_lo_hi_hi,header_lo_hi_lo,3'h0}; // @[Cat.scala 30:58]
  wire [1:0] _isLastState_T = a_hasData ? 2'h3 : 2'h2; // @[SinkA.scala 59:34]
  wire  isLastState = state == _isLastState_T; // @[SinkA.scala 59:27]
  wire [31:0] _io_q_bits_data_WIRE_1 = inject_io_o_bits_address; // @[SinkA.scala 63:25 SinkA.scala 63:25]
  wire [31:0] _GEN_39 = 2'h1 == state ? _io_q_bits_data_WIRE_1 : header; // @[SinkA.scala 63:19 SinkA.scala 63:19]
  wire [31:0] _GEN_40 = 2'h2 == state ? 32'h0 : _GEN_39; // @[SinkA.scala 63:19 SinkA.scala 63:19]
  wire [31:0] _io_q_bits_data_WIRE_3 = inject_io_o_bits_data; // @[SinkA.scala 63:25 SinkA.scala 63:25]
  wire [2:0] io_q_bits_beats_shiftAmount = header_hi_lo[2:0]; // @[OneHot.scala 64:49]
  wire [7:0] _io_q_bits_beats_T_1 = 8'h1 << io_q_bits_beats_shiftAmount; // @[OneHot.scala 65:12]
  wire [3:0] io_q_bits_beats_hi = _io_q_bits_beats_T_1[6:3]; // @[Parameters.scala 102:62]
  wire  io_q_bits_beats_lo = inject_io_o_bits_size <= 3'h2; // @[Parameters.scala 102:83]
  wire [4:0] _io_q_bits_beats_T_3 = {io_q_bits_beats_hi,io_q_bits_beats_lo}; // @[Cat.scala 30:58]
  wire [4:0] _io_q_bits_beats_T_4 = a_hasData ? _io_q_bits_beats_T_3 : 5'h0; // @[SinkA.scala 64:25]
  wire [4:0] _io_q_bits_beats_T_6 = _io_q_bits_beats_T_4 + 5'h3; // @[SinkA.scala 64:76]
  wire  io_q_bits_beats_hi_1 = _io_q_bits_beats_T_1[6]; // @[Parameters.scala 107:62]
  wire  io_q_bits_beats_lo_1 = inject_io_o_bits_size <= 3'h5; // @[Parameters.scala 107:83]
  wire [1:0] _io_q_bits_beats_T_10 = {io_q_bits_beats_hi_1,io_q_bits_beats_lo_1}; // @[Cat.scala 30:58]
  wire [1:0] _io_q_bits_beats_T_11 = a_partial ? _io_q_bits_beats_T_10 : 2'h0; // @[SinkA.scala 65:25]
  wire [4:0] _GEN_42 = {{3'd0}, _io_q_bits_beats_T_11}; // @[SinkA.scala 64:86]
  wire [4:0] _io_q_bits_beats_T_13 = _io_q_bits_beats_T_6 + _GEN_42; // @[SinkA.scala 64:86]
  PartialInjector inject ( // @[SinkA.scala 21:22]
    .clock(inject_clock),
    .reset(inject_reset),
    .io_i_last(inject_io_i_last),
    .io_o_last(inject_io_o_last),
    .io_i_ready(inject_io_i_ready),
    .io_i_valid(inject_io_i_valid),
    .io_i_bits_opcode(inject_io_i_bits_opcode),
    .io_i_bits_param(inject_io_i_bits_param),
    .io_i_bits_size(inject_io_i_bits_size),
    .io_i_bits_source(inject_io_i_bits_source),
    .io_i_bits_address(inject_io_i_bits_address),
    .io_i_bits_mask(inject_io_i_bits_mask),
    .io_i_bits_data(inject_io_i_bits_data),
    .io_o_ready(inject_io_o_ready),
    .io_o_valid(inject_io_o_valid),
    .io_o_bits_opcode(inject_io_o_bits_opcode),
    .io_o_bits_param(inject_io_o_bits_param),
    .io_o_bits_size(inject_io_o_bits_size),
    .io_o_bits_source(inject_io_o_bits_source),
    .io_o_bits_address(inject_io_o_bits_address),
    .io_o_bits_data(inject_io_o_bits_data)
  );
  Queue_2 inject_io_i_q ( // @[Decoupled.scala 296:21]
    .clock(inject_io_i_q_clock),
    .reset(inject_io_i_q_reset),
    .io_enq_ready(inject_io_i_q_io_enq_ready),
    .io_enq_valid(inject_io_i_q_io_enq_valid),
    .io_enq_bits_opcode(inject_io_i_q_io_enq_bits_opcode),
    .io_enq_bits_size(inject_io_i_q_io_enq_bits_size),
    .io_enq_bits_source(inject_io_i_q_io_enq_bits_source),
    .io_enq_bits_address(inject_io_i_q_io_enq_bits_address),
    .io_enq_bits_mask(inject_io_i_q_io_enq_bits_mask),
    .io_enq_bits_data(inject_io_i_q_io_enq_bits_data),
    .io_deq_ready(inject_io_i_q_io_deq_ready),
    .io_deq_valid(inject_io_i_q_io_deq_valid),
    .io_deq_bits_opcode(inject_io_i_q_io_deq_bits_opcode),
    .io_deq_bits_param(inject_io_i_q_io_deq_bits_param),
    .io_deq_bits_size(inject_io_i_q_io_deq_bits_size),
    .io_deq_bits_source(inject_io_i_q_io_deq_bits_source),
    .io_deq_bits_address(inject_io_i_q_io_deq_bits_address),
    .io_deq_bits_mask(inject_io_i_q_io_deq_bits_mask),
    .io_deq_bits_data(inject_io_i_q_io_deq_bits_data)
  );
  assign io_a_ready = inject_io_i_q_io_enq_ready; // @[Decoupled.scala 299:17]
  assign io_q_valid = inject_io_o_valid; // @[SinkA.scala 61:14]
  assign io_q_bits_data = 2'h3 == state ? _io_q_bits_data_WIRE_3 : _GEN_40; // @[SinkA.scala 63:19 SinkA.scala 63:19]
  assign io_q_bits_last = inject_io_o_last & isLastState; // @[SinkA.scala 62:29]
  assign io_q_bits_beats = {{2'd0}, _io_q_bits_beats_T_13}; // @[SinkA.scala 64:86]
  assign inject_clock = clock;
  assign inject_reset = reset;
  assign inject_io_i_last = inject_io_i_last_counter == 4'h1 | inject_io_i_last_beats1 == 4'h0; // @[Edges.scala 231:37]
  assign inject_io_i_valid = inject_io_i_q_io_deq_valid; // @[SinkA.scala 22:15]
  assign inject_io_i_bits_opcode = inject_io_i_q_io_deq_bits_opcode; // @[SinkA.scala 22:15]
  assign inject_io_i_bits_param = inject_io_i_q_io_deq_bits_param; // @[SinkA.scala 22:15]
  assign inject_io_i_bits_size = inject_io_i_q_io_deq_bits_size; // @[SinkA.scala 22:15]
  assign inject_io_i_bits_source = inject_io_i_q_io_deq_bits_source; // @[SinkA.scala 22:15]
  assign inject_io_i_bits_address = inject_io_i_q_io_deq_bits_address; // @[SinkA.scala 22:15]
  assign inject_io_i_bits_mask = inject_io_i_q_io_deq_bits_mask; // @[SinkA.scala 22:15]
  assign inject_io_i_bits_data = inject_io_i_q_io_deq_bits_data; // @[SinkA.scala 22:15]
  assign inject_io_o_ready = io_q_ready & isLastState; // @[SinkA.scala 60:25]
  assign inject_io_i_q_clock = clock;
  assign inject_io_i_q_reset = reset;
  assign inject_io_i_q_io_enq_valid = io_a_valid; // @[Decoupled.scala 297:22]
  assign inject_io_i_q_io_enq_bits_opcode = io_a_bits_opcode; // @[Decoupled.scala 298:21]
  assign inject_io_i_q_io_enq_bits_size = io_a_bits_size; // @[Decoupled.scala 298:21]
  assign inject_io_i_q_io_enq_bits_source = io_a_bits_source; // @[Decoupled.scala 298:21]
  assign inject_io_i_q_io_enq_bits_address = io_a_bits_address; // @[Decoupled.scala 298:21]
  assign inject_io_i_q_io_enq_bits_mask = io_a_bits_mask; // @[Decoupled.scala 298:21]
  assign inject_io_i_q_io_enq_bits_data = io_a_bits_data; // @[Decoupled.scala 298:21]
  assign inject_io_i_q_io_deq_ready = inject_io_i_ready; // @[SinkA.scala 22:15]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      inject_io_i_last_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_inject_io_i_last_T) begin // @[Edges.scala 234:17]
      if (inject_io_i_last_first) begin // @[Edges.scala 235:21]
        if (inject_io_i_last_beats1_opdata) begin // @[Edges.scala 220:14]
          inject_io_i_last_counter <= inject_io_i_last_beats1_decode;
        end else begin
          inject_io_i_last_counter <= 4'h0;
        end
      end else begin
        inject_io_i_last_counter <= inject_io_i_last_counter1;
      end
    end
    if (reset) begin // @[SinkA.scala 30:22]
      state <= 2'h0; // @[SinkA.scala 30:22]
    end else if (_T) begin // @[SinkA.scala 36:22]
      if (_T_1) begin // @[Conditional.scala 40:58]
        state <= 2'h1; // @[SinkA.scala 38:31]
      end else if (_T_2) begin // @[Conditional.scala 39:67]
        state <= 2'h2; // @[SinkA.scala 39:31]
      end else begin
        state <= _GEN_2;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inject_io_i_last_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinkB(
  input         clock,
  input         reset,
  input         io_q_ready,
  output        io_q_valid,
  output [31:0] io_q_bits_data,
  output        io_q_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[SinkB.scala 25:22]
  wire  _T = io_q_ready & io_q_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_1 = _T_4 ? 2'h0 : state; // @[Conditional.scala 39:67 SinkB.scala 36:31 SinkB.scala 25:22]
  wire [1:0] _GEN_2 = _T_3 ? 2'h0 : _GEN_1; // @[Conditional.scala 39:67 SinkB.scala 35:31]
  wire [31:0] _GEN_7 = 2'h1 == state ? 32'h0 : 32'h1; // @[SinkB.scala 60:19 SinkB.scala 60:19]
  wire [31:0] _GEN_8 = 2'h2 == state ? 32'h0 : _GEN_7; // @[SinkB.scala 60:19 SinkB.scala 60:19]
  assign io_q_valid = 1'h0; // @[SinkB.scala 58:14]
  assign io_q_bits_data = 2'h3 == state ? 32'h0 : _GEN_8; // @[SinkB.scala 60:19 SinkB.scala 60:19]
  assign io_q_bits_last = state == 2'h2; // @[SinkB.scala 56:27]
  always @(posedge clock) begin
    if (reset) begin // @[SinkB.scala 25:22]
      state <= 2'h0; // @[SinkB.scala 25:22]
    end else if (_T) begin // @[SinkB.scala 31:22]
      if (_T_1) begin // @[Conditional.scala 40:58]
        state <= 2'h1; // @[SinkB.scala 33:31]
      end else if (_T_2) begin // @[Conditional.scala 39:67]
        state <= 2'h2; // @[SinkB.scala 34:31]
      end else begin
        state <= _GEN_2;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinkC(
  input         clock,
  input         reset,
  input         io_q_ready,
  output        io_q_valid,
  output [31:0] io_q_bits_data,
  output        io_q_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[SinkC.scala 27:22]
  wire  _T = io_q_ready & io_q_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_1 = _T_4 ? 2'h0 : state; // @[Conditional.scala 39:67 SinkC.scala 38:31 SinkC.scala 27:22]
  wire [1:0] _GEN_2 = _T_3 ? 2'h0 : _GEN_1; // @[Conditional.scala 39:67 SinkC.scala 37:31]
  wire [31:0] _GEN_39 = 2'h1 == state ? 32'h0 : 32'h2; // @[SinkC.scala 62:19 SinkC.scala 62:19]
  wire [31:0] _GEN_40 = 2'h2 == state ? 32'h0 : _GEN_39; // @[SinkC.scala 62:19 SinkC.scala 62:19]
  assign io_q_valid = 1'h0; // @[SinkC.scala 60:14]
  assign io_q_bits_data = 2'h3 == state ? 32'h0 : _GEN_40; // @[SinkC.scala 62:19 SinkC.scala 62:19]
  assign io_q_bits_last = state == 2'h2; // @[SinkC.scala 58:27]
  always @(posedge clock) begin
    if (reset) begin // @[SinkC.scala 27:22]
      state <= 2'h0; // @[SinkC.scala 27:22]
    end else if (_T) begin // @[SinkC.scala 33:22]
      if (_T_1) begin // @[Conditional.scala 40:58]
        state <= 2'h1; // @[SinkC.scala 35:31]
      end else if (_T_2) begin // @[Conditional.scala 39:67]
        state <= 2'h2; // @[SinkC.scala 36:31]
      end else begin
        state <= _GEN_2;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_5(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [5:0]  io_enq_bits_source,
  input         io_enq_bits_denied,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [5:0]  io_deq_bits_source,
  output        io_deq_bits_sink,
  output        io_deq_bits_denied,
  output [31:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_param [0:0]; // @[Decoupled.scala 218:16]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [5:0] ram_source [0:0]; // @[Decoupled.scala 218:16]
  wire [5:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [5:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_sink [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sink_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_denied [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_data [0:0]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_14 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 249:27 Decoupled.scala 249:36]
  wire  do_enq = empty ? _GEN_14 : _do_enq_T; // @[Decoupled.scala 246:18]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 246:18 Decoupled.scala 248:14]
  assign ram_opcode_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = 1'h0;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_param_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = 1'h0;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = 1'h0;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_sink_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_sink_MPORT_data = 1'h0;
  assign ram_sink_MPORT_addr = 1'h0;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_denied_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = 1'h0;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_14 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 245:25 Decoupled.scala 245:40 Decoupled.scala 240:16]
  assign io_deq_bits_opcode = empty ? io_enq_bits_opcode : ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_param = empty ? io_enq_bits_param : ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_source = empty ? io_enq_bits_source : ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_sink = empty ? 1'h0 : ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_denied = empty ? io_enq_bits_denied : ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      if (empty) begin // @[Decoupled.scala 246:18]
        if (io_deq_ready) begin // @[Decoupled.scala 249:27]
          maybe_full <= 1'h0; // @[Decoupled.scala 249:36]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinkD(
  input         clock,
  input         reset,
  output        io_d_ready,
  input         io_d_valid,
  input  [2:0]  io_d_bits_opcode,
  input  [1:0]  io_d_bits_param,
  input  [2:0]  io_d_bits_size,
  input  [5:0]  io_d_bits_source,
  input         io_d_bits_denied,
  input  [31:0] io_d_bits_data,
  input         io_q_ready,
  output        io_q_valid,
  output [31:0] io_q_bits_data,
  output        io_q_bits_last,
  output [6:0]  io_q_bits_beats,
  output        io_a_tlSource_valid,
  output [5:0]  io_a_tlSource_bits,
  input  [15:0] io_a_clSource,
  output        io_c_tlSource_valid,
  output [5:0]  io_c_tlSource_bits,
  input  [15:0] io_c_clSource
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  d_clock; // @[Decoupled.scala 296:21]
  wire  d_reset; // @[Decoupled.scala 296:21]
  wire  d_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  d_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] d_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [1:0] d_io_enq_bits_param; // @[Decoupled.scala 296:21]
  wire [2:0] d_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [5:0] d_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire  d_io_enq_bits_denied; // @[Decoupled.scala 296:21]
  wire [31:0] d_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  d_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  d_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] d_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [1:0] d_io_deq_bits_param; // @[Decoupled.scala 296:21]
  wire [2:0] d_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [5:0] d_io_deq_bits_source; // @[Decoupled.scala 296:21]
  wire  d_io_deq_bits_sink; // @[Decoupled.scala 296:21]
  wire  d_io_deq_bits_denied; // @[Decoupled.scala 296:21]
  wire [31:0] d_io_deq_bits_data; // @[Decoupled.scala 296:21]
  reg [1:0] state; // @[SinkD.scala 20:22]
  wire  _d_last_T = d_io_deq_ready & d_io_deq_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_last_beats1_decode_T_1 = 13'h3f << d_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_last_beats1_decode_T_3 = ~_d_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_last_beats1_decode = _d_last_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_last_beats1_opdata = d_io_deq_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [3:0] d_last_beats1 = d_last_beats1_opdata ? d_last_beats1_decode : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] d_last_counter; // @[Edges.scala 228:27]
  wire [3:0] d_last_counter1 = d_last_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_last_first = d_last_counter == 4'h0; // @[Edges.scala 230:25]
  wire  d_last = d_last_counter == 4'h1 | d_last_beats1 == 4'h0; // @[Edges.scala 231:37]
  wire  d_grant = d_io_deq_bits_opcode == 3'h4 | d_io_deq_bits_opcode == 3'h5; // @[SinkD.scala 29:52]
  wire  _T = io_q_ready & io_q_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T = d_last_beats1_opdata ? 2'h2 : 2'h0; // @[SinkD.scala 33:58]
  wire  _T_2 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T_3 = d_last ? 2'h0 : 2'h2; // @[SinkD.scala 35:37]
  wire [1:0] _GEN_1 = _T_3 ? _state_T_3 : state; // @[Conditional.scala 39:67 SinkD.scala 35:31 SinkD.scala 20:22]
  wire  relack = d_io_deq_bits_opcode == 3'h6; // @[SinkD.scala 40:30]
  wire  _io_a_tlSource_valid_T_2 = _T & state == 2'h0; // @[SinkD.scala 41:38]
  wire [2:0] header_hi_hi_lo = d_io_deq_bits_source[5:3]; // @[SinkD.scala 52:28]
  wire [15:0] header_hi_hi_hi = relack ? io_c_clSource : io_a_clSource; // @[SinkD.scala 53:17]
  wire [3:0] header_hi_lo = {{1'd0}, d_io_deq_bits_size}; // @[Parameters.scala 80:35]
  wire [2:0] header_lo_hi_lo = d_io_deq_bits_opcode; // @[Parameters.scala 80:35]
  wire [31:0] header = {header_hi_hi_hi,header_hi_hi_lo,header_hi_lo,d_io_deq_bits_denied,d_io_deq_bits_param,
    header_lo_hi_lo,3'h3}; // @[Cat.scala 30:58]
  wire [1:0] _isLastState_T = d_grant ? 2'h1 : 2'h0; // @[SinkD.scala 55:57]
  wire [1:0] _isLastState_T_1 = d_last_beats1_opdata ? 2'h2 : _isLastState_T; // @[SinkD.scala 55:34]
  wire  isLastState = state == _isLastState_T_1; // @[SinkD.scala 55:27]
  wire [31:0] _io_q_bits_data_WIRE_1 = {{31'd0}, d_io_deq_bits_sink}; // @[SinkD.scala 59:25 SinkD.scala 59:25]
  wire [31:0] _GEN_6 = 2'h1 == state ? _io_q_bits_data_WIRE_1 : header; // @[SinkD.scala 59:19 SinkD.scala 59:19]
  wire [31:0] _io_q_bits_data_WIRE_2 = d_io_deq_bits_data; // @[SinkD.scala 59:25 SinkD.scala 59:25]
  wire [2:0] io_q_bits_beats_shiftAmount = header_hi_lo[2:0]; // @[OneHot.scala 64:49]
  wire [7:0] _io_q_bits_beats_T_1 = 8'h1 << io_q_bits_beats_shiftAmount; // @[OneHot.scala 65:12]
  wire [3:0] io_q_bits_beats_hi = _io_q_bits_beats_T_1[6:3]; // @[Parameters.scala 102:62]
  wire  io_q_bits_beats_lo = d_io_deq_bits_size <= 3'h2; // @[Parameters.scala 102:83]
  wire [4:0] _io_q_bits_beats_T_3 = {io_q_bits_beats_hi,io_q_bits_beats_lo}; // @[Cat.scala 30:58]
  wire [4:0] _io_q_bits_beats_T_4 = d_last_beats1_opdata ? _io_q_bits_beats_T_3 : 5'h0; // @[SinkD.scala 60:25]
  wire [4:0] _io_q_bits_beats_T_6 = _io_q_bits_beats_T_4 + 5'h1; // @[SinkD.scala 60:76]
  wire [4:0] _GEN_8 = {{4'd0}, d_grant}; // @[SinkD.scala 60:86]
  wire [4:0] _io_q_bits_beats_T_8 = _io_q_bits_beats_T_6 + _GEN_8; // @[SinkD.scala 60:86]
  Queue_5 d ( // @[Decoupled.scala 296:21]
    .clock(d_clock),
    .reset(d_reset),
    .io_enq_ready(d_io_enq_ready),
    .io_enq_valid(d_io_enq_valid),
    .io_enq_bits_opcode(d_io_enq_bits_opcode),
    .io_enq_bits_param(d_io_enq_bits_param),
    .io_enq_bits_size(d_io_enq_bits_size),
    .io_enq_bits_source(d_io_enq_bits_source),
    .io_enq_bits_denied(d_io_enq_bits_denied),
    .io_enq_bits_data(d_io_enq_bits_data),
    .io_deq_ready(d_io_deq_ready),
    .io_deq_valid(d_io_deq_valid),
    .io_deq_bits_opcode(d_io_deq_bits_opcode),
    .io_deq_bits_param(d_io_deq_bits_param),
    .io_deq_bits_size(d_io_deq_bits_size),
    .io_deq_bits_source(d_io_deq_bits_source),
    .io_deq_bits_sink(d_io_deq_bits_sink),
    .io_deq_bits_denied(d_io_deq_bits_denied),
    .io_deq_bits_data(d_io_deq_bits_data)
  );
  assign io_d_ready = d_io_enq_ready; // @[Decoupled.scala 299:17]
  assign io_q_valid = d_io_deq_valid; // @[SinkD.scala 57:14]
  assign io_q_bits_data = 2'h2 == state ? _io_q_bits_data_WIRE_2 : _GEN_6; // @[SinkD.scala 59:19 SinkD.scala 59:19]
  assign io_q_bits_last = d_last & isLastState; // @[SinkD.scala 58:29]
  assign io_q_bits_beats = {{2'd0}, _io_q_bits_beats_T_8}; // @[SinkD.scala 60:86]
  assign io_a_tlSource_valid = _T & state == 2'h0 & ~relack; // @[SinkD.scala 41:60]
  assign io_a_tlSource_bits = d_io_deq_bits_source; // @[SinkD.scala 42:22]
  assign io_c_tlSource_valid = _io_a_tlSource_valid_T_2 & relack; // @[SinkD.scala 43:60]
  assign io_c_tlSource_bits = d_io_deq_bits_source; // @[SinkD.scala 44:22]
  assign d_clock = clock;
  assign d_reset = reset;
  assign d_io_enq_valid = io_d_valid; // @[Decoupled.scala 297:22]
  assign d_io_enq_bits_opcode = io_d_bits_opcode; // @[Decoupled.scala 298:21]
  assign d_io_enq_bits_param = io_d_bits_param; // @[Decoupled.scala 298:21]
  assign d_io_enq_bits_size = io_d_bits_size; // @[Decoupled.scala 298:21]
  assign d_io_enq_bits_source = io_d_bits_source; // @[Decoupled.scala 298:21]
  assign d_io_enq_bits_denied = io_d_bits_denied; // @[Decoupled.scala 298:21]
  assign d_io_enq_bits_data = io_d_bits_data; // @[Decoupled.scala 298:21]
  assign d_io_deq_ready = io_q_ready & isLastState; // @[SinkD.scala 56:25]
  always @(posedge clock) begin
    if (reset) begin // @[SinkD.scala 20:22]
      state <= 2'h0; // @[SinkD.scala 20:22]
    end else if (_T) begin // @[SinkD.scala 31:22]
      if (_T_1) begin // @[Conditional.scala 40:58]
        if (d_grant) begin // @[SinkD.scala 33:37]
          state <= 2'h1;
        end else begin
          state <= _state_T;
        end
      end else if (_T_2) begin // @[Conditional.scala 39:67]
        state <= _state_T; // @[SinkD.scala 34:31]
      end else begin
        state <= _GEN_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_last_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_last_T) begin // @[Edges.scala 234:17]
      if (d_last_first) begin // @[Edges.scala 235:21]
        if (d_last_beats1_opdata) begin // @[Edges.scala 220:14]
          d_last_counter <= d_last_beats1_decode;
        end else begin
          d_last_counter <= 4'h0;
        end
      end else begin
        d_last_counter <= d_last_counter1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  d_last_counter = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinkE(
  output [31:0] io_q_bits_data,
  input  [15:0] io_d_clSink
);
  wire [22:0] header_hi = {io_d_clSink,3'h0,4'h0}; // @[Cat.scala 30:58]
  assign io_q_bits_data = {header_hi,9'h4}; // @[Cat.scala 30:58]
endmodule
module CAM(
  input         clock,
  input         reset,
  output        io_alloc_ready,
  input         io_alloc_valid,
  input  [15:0] io_alloc_bits,
  output [2:0]  io_key,
  input         io_free_valid,
  input  [2:0]  io_free_bits,
  output [15:0] io_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] data [0:7]; // @[CAM.scala 22:17]
  wire [15:0] data_io_data_MPORT_data; // @[CAM.scala 22:17]
  wire [2:0] data_io_data_MPORT_addr; // @[CAM.scala 22:17]
  wire [15:0] data_MPORT_data; // @[CAM.scala 22:17]
  wire [2:0] data_MPORT_addr; // @[CAM.scala 22:17]
  wire  data_MPORT_mask; // @[CAM.scala 22:17]
  wire  data_MPORT_en; // @[CAM.scala 22:17]
  reg [7:0] free; // @[CAM.scala 21:21]
  wire [8:0] _free_sel_T = {free, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _free_sel_T_2 = free | _free_sel_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _free_sel_T_3 = {_free_sel_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _free_sel_T_5 = _free_sel_T_2 | _free_sel_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _free_sel_T_6 = {_free_sel_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _free_sel_T_8 = _free_sel_T_5 | _free_sel_T_6[7:0]; // @[package.scala 244:43]
  wire [8:0] _free_sel_T_10 = {_free_sel_T_8, 1'h0}; // @[CAM.scala 24:39]
  wire [8:0] _free_sel_T_11 = ~_free_sel_T_10; // @[CAM.scala 24:18]
  wire [8:0] _GEN_5 = {{1'd0}, free}; // @[CAM.scala 24:45]
  wire [8:0] free_sel = _free_sel_T_11 & _GEN_5; // @[CAM.scala 24:45]
  wire [3:0] io_key_hi = free_sel[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] io_key_lo = free_sel[3:0]; // @[OneHot.scala 31:18]
  wire  io_key_hi_1 = |io_key_hi; // @[OneHot.scala 32:14]
  wire [3:0] _io_key_T = io_key_hi | io_key_lo; // @[OneHot.scala 32:28]
  wire [1:0] io_key_hi_2 = _io_key_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_key_lo_1 = _io_key_T[1:0]; // @[OneHot.scala 31:18]
  wire  io_key_hi_3 = |io_key_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _io_key_T_1 = io_key_hi_2 | io_key_lo_1; // @[OneHot.scala 32:28]
  wire  io_key_lo_2 = _io_key_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] io_key_lo_3 = {io_key_hi_3,io_key_lo_2}; // @[Cat.scala 30:58]
  wire  _T = io_alloc_ready & io_alloc_valid; // @[Decoupled.scala 40:37]
  wire  bypass = _T & io_free_bits == io_key; // @[CAM.scala 31:32]
  wire [8:0] clr = _T ? free_sel : 9'h0; // @[CAM.scala 35:16]
  wire [7:0] _set_T = 8'h1 << io_free_bits; // @[OneHot.scala 58:35]
  wire [7:0] set = io_free_valid ? _set_T : 8'h0; // @[CAM.scala 36:16]
  wire [8:0] _free_T = ~clr; // @[CAM.scala 37:19]
  wire [8:0] _free_T_1 = _GEN_5 & _free_T; // @[CAM.scala 37:17]
  wire [8:0] _GEN_7 = {{1'd0}, set}; // @[CAM.scala 37:25]
  wire [8:0] _free_T_2 = _free_T_1 | _GEN_7; // @[CAM.scala 37:25]
  assign data_io_data_MPORT_addr = io_free_bits;
  assign data_io_data_MPORT_data = data[data_io_data_MPORT_addr]; // @[CAM.scala 22:17]
  assign data_MPORT_data = io_alloc_bits;
  assign data_MPORT_addr = io_key;
  assign data_MPORT_mask = 1'h1;
  assign data_MPORT_en = io_alloc_ready & io_alloc_valid;
  assign io_alloc_ready = |free; // @[CAM.scala 27:26]
  assign io_key = {io_key_hi_1,io_key_lo_3}; // @[Cat.scala 30:58]
  assign io_data = bypass ? io_alloc_bits : data_io_data_MPORT_data; // @[CAM.scala 32:17]
  always @(posedge clock) begin
    if(data_MPORT_en & data_MPORT_mask) begin
      data[data_MPORT_addr] <= data_MPORT_data; // @[CAM.scala 22:17]
    end
    if (reset) begin // @[CAM.scala 21:21]
      free <= 8'hff; // @[CAM.scala 21:21]
    end else begin
      free <= _free_T_2[7:0]; // @[CAM.scala 37:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  free = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ParitalExtractor(
  input         clock,
  input         reset,
  input         io_last,
  output        io_i_ready,
  input         io_i_valid,
  input  [2:0]  io_i_bits_opcode,
  input  [2:0]  io_i_bits_param,
  input  [2:0]  io_i_bits_size,
  input  [5:0]  io_i_bits_source,
  input  [31:0] io_i_bits_address,
  input  [3:0]  io_i_bits_mask,
  input  [31:0] io_i_bits_data,
  input         io_o_ready,
  output        io_o_valid,
  output [2:0]  io_o_bits_opcode,
  output [2:0]  io_o_bits_param,
  output [2:0]  io_o_bits_size,
  output [5:0]  io_o_bits_source,
  output [31:0] io_o_bits_address,
  output [3:0]  io_o_bits_mask,
  output [31:0] io_o_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] state; // @[Partial.scala 29:23]
  reg [31:0] shift; // @[Partial.scala 30:19]
  wire  enable = io_i_bits_opcode == 3'h1; // @[Partial.scala 31:25]
  wire  empty = state == 4'h0; // @[Partial.scala 32:22]
  wire [5:0] _wide_T = {state, 2'h0}; // @[Partial.scala 35:42]
  wire [94:0] _GEN_12 = {{63'd0}, io_i_bits_data}; // @[Partial.scala 35:32]
  wire [94:0] _wide_T_1 = _GEN_12 << _wide_T; // @[Partial.scala 35:32]
  wire [94:0] _GEN_13 = {{63'd0}, shift}; // @[Partial.scala 35:22]
  wire [94:0] wide = _GEN_13 | _wide_T_1; // @[Partial.scala 35:22]
  wire [31:0] _io_o_bits_data_T_4 = {wide[35:28],wide[26:19],wide[17:10],wide[8:1]}; // @[Partial.scala 36:64]
  wire [3:0] _io_o_bits_mask_T_4 = {wide[27],wide[18],wide[9],wide[0]}; // @[Partial.scala 37:51]
  wire  _GEN_0 = empty | io_o_ready; // @[Partial.scala 40:18 Partial.scala 41:18 Partial.scala 17:8]
  wire  _GEN_1 = empty ? 1'h0 : io_i_valid; // @[Partial.scala 40:18 Partial.scala 42:18 Partial.scala 17:8]
  wire  _T = io_i_ready & io_i_valid; // @[Decoupled.scala 40:37]
  wire [58:0] _shift_T_1 = empty ? {{27'd0}, io_i_bits_data} : wide[94:36]; // @[Partial.scala 47:19]
  wire [3:0] _state_T_1 = state - 4'h1; // @[Partial.scala 48:22]
  wire [3:0] _GEN_2 = empty ? 4'h8 : _state_T_1; // @[Partial.scala 49:22 Partial.scala 49:30 Partial.scala 48:13]
  wire [58:0] _GEN_4 = _T ? _shift_T_1 : {{27'd0}, shift}; // @[Partial.scala 46:24 Partial.scala 47:13 Partial.scala 30:19]
  wire [58:0] _GEN_10 = enable ? _GEN_4 : {{27'd0}, shift}; // @[Partial.scala 34:17 Partial.scala 30:19]
  assign io_i_ready = enable ? _GEN_0 : io_o_ready; // @[Partial.scala 34:17 Partial.scala 17:8]
  assign io_o_valid = enable ? _GEN_1 : io_i_valid; // @[Partial.scala 34:17 Partial.scala 17:8]
  assign io_o_bits_opcode = io_i_bits_opcode; // @[Partial.scala 17:8]
  assign io_o_bits_param = io_i_bits_param; // @[Partial.scala 17:8]
  assign io_o_bits_size = io_i_bits_size; // @[Partial.scala 17:8]
  assign io_o_bits_source = io_i_bits_source; // @[Partial.scala 17:8]
  assign io_o_bits_address = io_i_bits_address; // @[Partial.scala 17:8]
  assign io_o_bits_mask = enable ? _io_o_bits_mask_T_4 : io_i_bits_mask; // @[Partial.scala 34:17 Partial.scala 37:12 Partial.scala 17:8]
  assign io_o_bits_data = enable ? _io_o_bits_data_T_4 : io_i_bits_data; // @[Partial.scala 34:17 Partial.scala 36:12 Partial.scala 17:8]
  always @(posedge clock) begin
    if (reset) begin // @[Partial.scala 29:23]
      state <= 4'h0; // @[Partial.scala 29:23]
    end else if (enable) begin // @[Partial.scala 34:17]
      if (_T) begin // @[Partial.scala 46:24]
        if (io_last) begin // @[Partial.scala 50:22]
          state <= 4'h0; // @[Partial.scala 50:30]
        end else begin
          state <= _GEN_2;
        end
      end
    end
    shift <= _GEN_10[31:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  shift = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SourceA(
  input         clock,
  input         reset,
  input         io_a_ready,
  output        io_a_valid,
  output [2:0]  io_a_bits_opcode,
  output [2:0]  io_a_bits_param,
  output [2:0]  io_a_bits_size,
  output [5:0]  io_a_bits_source,
  output [31:0] io_a_bits_address,
  output [3:0]  io_a_bits_mask,
  output [31:0] io_a_bits_data,
  output        io_q_ready,
  input         io_q_valid,
  input  [31:0] io_q_bits,
  input         io_d_tlSource_valid,
  input  [5:0]  io_d_tlSource_bits,
  output [15:0] io_d_clSource
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  cams_0_clock; // @[SourceA.scala 21:11]
  wire  cams_0_reset; // @[SourceA.scala 21:11]
  wire  cams_0_io_alloc_ready; // @[SourceA.scala 21:11]
  wire  cams_0_io_alloc_valid; // @[SourceA.scala 21:11]
  wire [15:0] cams_0_io_alloc_bits; // @[SourceA.scala 21:11]
  wire [2:0] cams_0_io_key; // @[SourceA.scala 21:11]
  wire  cams_0_io_free_valid; // @[SourceA.scala 21:11]
  wire [2:0] cams_0_io_free_bits; // @[SourceA.scala 21:11]
  wire [15:0] cams_0_io_data; // @[SourceA.scala 21:11]
  wire  cams_1_clock; // @[SourceA.scala 21:11]
  wire  cams_1_reset; // @[SourceA.scala 21:11]
  wire  cams_1_io_alloc_ready; // @[SourceA.scala 21:11]
  wire  cams_1_io_alloc_valid; // @[SourceA.scala 21:11]
  wire [15:0] cams_1_io_alloc_bits; // @[SourceA.scala 21:11]
  wire [2:0] cams_1_io_key; // @[SourceA.scala 21:11]
  wire  cams_1_io_free_valid; // @[SourceA.scala 21:11]
  wire [2:0] cams_1_io_free_bits; // @[SourceA.scala 21:11]
  wire [15:0] cams_1_io_data; // @[SourceA.scala 21:11]
  wire  cams_2_clock; // @[SourceA.scala 21:11]
  wire  cams_2_reset; // @[SourceA.scala 21:11]
  wire  cams_2_io_alloc_ready; // @[SourceA.scala 21:11]
  wire  cams_2_io_alloc_valid; // @[SourceA.scala 21:11]
  wire [15:0] cams_2_io_alloc_bits; // @[SourceA.scala 21:11]
  wire [2:0] cams_2_io_key; // @[SourceA.scala 21:11]
  wire  cams_2_io_free_valid; // @[SourceA.scala 21:11]
  wire [2:0] cams_2_io_free_bits; // @[SourceA.scala 21:11]
  wire [15:0] cams_2_io_data; // @[SourceA.scala 21:11]
  wire  cams_3_clock; // @[SourceA.scala 21:11]
  wire  cams_3_reset; // @[SourceA.scala 21:11]
  wire  cams_3_io_alloc_ready; // @[SourceA.scala 21:11]
  wire  cams_3_io_alloc_valid; // @[SourceA.scala 21:11]
  wire [15:0] cams_3_io_alloc_bits; // @[SourceA.scala 21:11]
  wire [2:0] cams_3_io_key; // @[SourceA.scala 21:11]
  wire  cams_3_io_free_valid; // @[SourceA.scala 21:11]
  wire [2:0] cams_3_io_free_bits; // @[SourceA.scala 21:11]
  wire [15:0] cams_3_io_data; // @[SourceA.scala 21:11]
  wire  cams_4_clock; // @[SourceA.scala 21:11]
  wire  cams_4_reset; // @[SourceA.scala 21:11]
  wire  cams_4_io_alloc_ready; // @[SourceA.scala 21:11]
  wire  cams_4_io_alloc_valid; // @[SourceA.scala 21:11]
  wire [15:0] cams_4_io_alloc_bits; // @[SourceA.scala 21:11]
  wire [2:0] cams_4_io_key; // @[SourceA.scala 21:11]
  wire  cams_4_io_free_valid; // @[SourceA.scala 21:11]
  wire [2:0] cams_4_io_free_bits; // @[SourceA.scala 21:11]
  wire [15:0] cams_4_io_data; // @[SourceA.scala 21:11]
  wire  cams_5_clock; // @[SourceA.scala 21:11]
  wire  cams_5_reset; // @[SourceA.scala 21:11]
  wire  cams_5_io_alloc_ready; // @[SourceA.scala 21:11]
  wire  cams_5_io_alloc_valid; // @[SourceA.scala 21:11]
  wire [15:0] cams_5_io_alloc_bits; // @[SourceA.scala 21:11]
  wire [2:0] cams_5_io_key; // @[SourceA.scala 21:11]
  wire  cams_5_io_free_valid; // @[SourceA.scala 21:11]
  wire [2:0] cams_5_io_free_bits; // @[SourceA.scala 21:11]
  wire [15:0] cams_5_io_data; // @[SourceA.scala 21:11]
  wire  cams_6_clock; // @[SourceA.scala 21:11]
  wire  cams_6_reset; // @[SourceA.scala 21:11]
  wire  cams_6_io_alloc_ready; // @[SourceA.scala 21:11]
  wire  cams_6_io_alloc_valid; // @[SourceA.scala 21:11]
  wire [15:0] cams_6_io_alloc_bits; // @[SourceA.scala 21:11]
  wire [2:0] cams_6_io_key; // @[SourceA.scala 21:11]
  wire  cams_6_io_free_valid; // @[SourceA.scala 21:11]
  wire [2:0] cams_6_io_free_bits; // @[SourceA.scala 21:11]
  wire [15:0] cams_6_io_data; // @[SourceA.scala 21:11]
  wire  cams_7_clock; // @[SourceA.scala 21:11]
  wire  cams_7_reset; // @[SourceA.scala 21:11]
  wire  cams_7_io_alloc_ready; // @[SourceA.scala 21:11]
  wire  cams_7_io_alloc_valid; // @[SourceA.scala 21:11]
  wire [15:0] cams_7_io_alloc_bits; // @[SourceA.scala 21:11]
  wire [2:0] cams_7_io_key; // @[SourceA.scala 21:11]
  wire  cams_7_io_free_valid; // @[SourceA.scala 21:11]
  wire [2:0] cams_7_io_free_bits; // @[SourceA.scala 21:11]
  wire [15:0] cams_7_io_data; // @[SourceA.scala 21:11]
  wire  extract_clock; // @[SourceA.scala 75:23]
  wire  extract_reset; // @[SourceA.scala 75:23]
  wire  extract_io_last; // @[SourceA.scala 75:23]
  wire  extract_io_i_ready; // @[SourceA.scala 75:23]
  wire  extract_io_i_valid; // @[SourceA.scala 75:23]
  wire [2:0] extract_io_i_bits_opcode; // @[SourceA.scala 75:23]
  wire [2:0] extract_io_i_bits_param; // @[SourceA.scala 75:23]
  wire [2:0] extract_io_i_bits_size; // @[SourceA.scala 75:23]
  wire [5:0] extract_io_i_bits_source; // @[SourceA.scala 75:23]
  wire [31:0] extract_io_i_bits_address; // @[SourceA.scala 75:23]
  wire [3:0] extract_io_i_bits_mask; // @[SourceA.scala 75:23]
  wire [31:0] extract_io_i_bits_data; // @[SourceA.scala 75:23]
  wire  extract_io_o_ready; // @[SourceA.scala 75:23]
  wire  extract_io_o_valid; // @[SourceA.scala 75:23]
  wire [2:0] extract_io_o_bits_opcode; // @[SourceA.scala 75:23]
  wire [2:0] extract_io_o_bits_param; // @[SourceA.scala 75:23]
  wire [2:0] extract_io_o_bits_size; // @[SourceA.scala 75:23]
  wire [5:0] extract_io_o_bits_source; // @[SourceA.scala 75:23]
  wire [31:0] extract_io_o_bits_address; // @[SourceA.scala 75:23]
  wire [3:0] extract_io_o_bits_mask; // @[SourceA.scala 75:23]
  wire [31:0] extract_io_o_bits_data; // @[SourceA.scala 75:23]
  reg [1:0] state; // @[SourceA.scala 25:22]
  wire [2:0] opcode = io_q_bits[5:3]; // @[Parameters.scala 92:19]
  wire [2:0] param = io_q_bits[8:6]; // @[Parameters.scala 93:19]
  wire [3:0] size = io_q_bits[12:9]; // @[Parameters.scala 94:19]
  wire [2:0] domain = io_q_bits[15:13]; // @[Parameters.scala 95:19]
  wire [15:0] source = io_q_bits[31:16]; // @[Parameters.scala 96:19]
  wire  enable = state == 2'h0; // @[SourceA.scala 32:24]
  reg [2:0] r_1; // @[Reg.scala 15:16]
  wire [2:0] _GEN_1 = enable ? opcode : r_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [2:0] r_2; // @[Reg.scala 15:16]
  reg [3:0] r_3; // @[Reg.scala 15:16]
  wire [3:0] _GEN_3 = enable ? size : r_3; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [2:0] r_4; // @[Reg.scala 15:16]
  wire [2:0] _GEN_4 = enable ? domain : r_4; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [15:0] r_5; // @[Reg.scala 15:16]
  wire  q_address0_enable = state == 2'h1; // @[SourceA.scala 32:24]
  reg [31:0] q_address0_r; // @[Reg.scala 15:16]
  wire [31:0] _GEN_6 = q_address0_enable ? io_q_bits : q_address0_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire  q_address1_enable = state == 2'h2; // @[SourceA.scala 32:24]
  reg [31:0] q_address1_r; // @[Reg.scala 15:16]
  wire [31:0] _GEN_7 = q_address1_enable ? io_q_bits : q_address1_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [4:0] q_last_count; // @[Parameters.scala 126:24]
  wire [2:0] q_last_beats_beats_shiftAmount = size[2:0]; // @[OneHot.scala 64:49]
  wire [7:0] _q_last_beats_beats_T_1 = 8'h1 << q_last_beats_beats_shiftAmount; // @[OneHot.scala 65:12]
  wire [3:0] q_last_beats_beats_hi = _q_last_beats_beats_T_1[6:3]; // @[Parameters.scala 102:62]
  wire  q_last_beats_beats_lo = size <= 4'h2; // @[Parameters.scala 102:83]
  wire [4:0] q_last_beats_beats = {q_last_beats_beats_hi,q_last_beats_beats_lo}; // @[Cat.scala 30:58]
  wire  q_last_beats_masks_hi = _q_last_beats_beats_T_1[6]; // @[Parameters.scala 107:62]
  wire  q_last_beats_masks_lo = size <= 4'h5; // @[Parameters.scala 107:83]
  wire [1:0] q_last_beats_masks = {q_last_beats_masks_hi,q_last_beats_masks_lo}; // @[Cat.scala 30:58]
  wire  q_last_beats_partial = opcode == 3'h1; // @[Parameters.scala 115:26]
  wire [4:0] _q_last_beats_a_T_1 = opcode[2] ? 5'h0 : q_last_beats_beats; // @[Parameters.scala 116:16]
  wire [4:0] _q_last_beats_a_T_3 = _q_last_beats_a_T_1 + 5'h2; // @[Parameters.scala 116:44]
  wire [1:0] _q_last_beats_a_T_4 = q_last_beats_partial ? q_last_beats_masks : 2'h0; // @[Parameters.scala 116:59]
  wire [4:0] _GEN_40 = {{3'd0}, _q_last_beats_a_T_4}; // @[Parameters.scala 116:54]
  wire [4:0] q_last_beats_a = _q_last_beats_a_T_3 + _GEN_40; // @[Parameters.scala 116:54]
  wire  q_last_first = q_last_count == 5'h0; // @[Parameters.scala 128:23]
  wire  q_last = q_last_count == 5'h1 | q_last_first & q_last_beats_a == 5'h0; // @[Parameters.scala 129:35]
  wire  _q_last_T = io_q_ready & io_q_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _q_last_count_T_1 = q_last_count - 5'h1; // @[Parameters.scala 130:56]
  wire  q_hasData = ~_GEN_1[2]; // @[SourceA.scala 45:19]
  wire  _a_first_T = state != 2'h3; // @[SourceA.scala 46:33]
  reg  a_first; // @[Reg.scala 15:16]
  wire  _T_2 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T = q_hasData ? 2'h3 : 2'h0; // @[SourceA.scala 52:37]
  wire  _T_5 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T_2 = ~q_last ? 2'h3 : 2'h0; // @[SourceA.scala 53:37]
  wire [1:0] _GEN_10 = _T_5 ? _state_T_2 : state; // @[Conditional.scala 39:67 SourceA.scala 53:31 SourceA.scala 25:22]
  wire [1:0] _GEN_11 = _T_4 ? _state_T : _GEN_10; // @[Conditional.scala 39:67 SourceA.scala 52:31]
  wire [63:0] q_address = {_GEN_7,_GEN_6}; // @[Cat.scala 30:58]
  wire  q_acq = _GEN_1 == 3'h6 | _GEN_1 == 3'h7; // @[SourceA.scala 59:52]
  wire [63:0] _exists_T = q_address ^ 64'h10000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_1 = {1'b0,$signed(_exists_T)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_3 = $signed(_exists_T_1) & -65'sh10000000; // @[Parameters.scala 137:52]
  wire  _exists_T_4 = $signed(_exists_T_3) == 65'sh0; // @[Parameters.scala 137:67]
  wire [63:0] _exists_T_5 = q_address ^ 64'h20000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_6 = {1'b0,$signed(_exists_T_5)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_8 = $signed(_exists_T_6) & -65'sh20000000; // @[Parameters.scala 137:52]
  wire  _exists_T_9 = $signed(_exists_T_8) == 65'sh0; // @[Parameters.scala 137:67]
  wire [63:0] _exists_T_10 = q_address ^ 64'h40000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_11 = {1'b0,$signed(_exists_T_10)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_13 = $signed(_exists_T_11) & -65'sh40000000; // @[Parameters.scala 137:52]
  wire  _exists_T_14 = $signed(_exists_T_13) == 65'sh0; // @[Parameters.scala 137:67]
  wire [63:0] _exists_T_15 = q_address ^ 64'h80000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_16 = {1'b0,$signed(_exists_T_15)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_18 = $signed(_exists_T_16) & -65'sh40000000; // @[Parameters.scala 137:52]
  wire  _exists_T_19 = $signed(_exists_T_18) == 65'sh0; // @[Parameters.scala 137:67]
  wire [63:0] _exists_T_20 = q_address ^ 64'hc0000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_21 = {1'b0,$signed(_exists_T_20)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_23 = $signed(_exists_T_21) & -65'sh20000000; // @[Parameters.scala 137:52]
  wire  _exists_T_24 = $signed(_exists_T_23) == 65'sh0; // @[Parameters.scala 137:67]
  wire  _exists_T_28 = _exists_T_4 | _exists_T_9 | _exists_T_14 | _exists_T_19 | _exists_T_24; // @[Parameters.scala 598:92]
  wire [63:0] _exists_T_29 = q_address ^ 64'h1000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_30 = {1'b0,$signed(_exists_T_29)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_32 = $signed(_exists_T_30) & -65'sh1000; // @[Parameters.scala 137:52]
  wire  _exists_T_33 = $signed(_exists_T_32) == 65'sh0; // @[Parameters.scala 137:67]
  wire  exists = _exists_T_28 | _exists_T_33; // @[Parameters.scala 622:64]
  wire [64:0] _writeOk_T_1 = {1'b0,$signed(q_address)}; // @[Parameters.scala 137:49]
  wire [64:0] _acquireOk_T_32 = $signed(_writeOk_T_1) & 65'shf0000000; // @[Parameters.scala 137:52]
  wire  acquireOk = $signed(_acquireOk_T_32) == 65'sh0; // @[Parameters.scala 137:67]
  wire  q_legal = exists & (~q_acq | acquireOk); // @[SourceA.scala 67:49]
  reg [2:0] source_r; // @[Reg.scala 15:16]
  wire [2:0] _source_WIRE_0 = cams_0_io_key; // @[SourceA.scala 71:22 SourceA.scala 71:22]
  wire [2:0] _source_WIRE_1 = cams_1_io_key; // @[SourceA.scala 71:22 SourceA.scala 71:22]
  wire [2:0] _GEN_16 = 3'h1 == _GEN_4 ? _source_WIRE_1 : _source_WIRE_0; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire [2:0] _source_WIRE_2 = cams_2_io_key; // @[SourceA.scala 71:22 SourceA.scala 71:22]
  wire [2:0] _GEN_17 = 3'h2 == _GEN_4 ? _source_WIRE_2 : _GEN_16; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire [2:0] _source_WIRE_3 = cams_3_io_key; // @[SourceA.scala 71:22 SourceA.scala 71:22]
  wire [2:0] _GEN_18 = 3'h3 == _GEN_4 ? _source_WIRE_3 : _GEN_17; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire [2:0] _source_WIRE_4 = cams_4_io_key; // @[SourceA.scala 71:22 SourceA.scala 71:22]
  wire [2:0] _GEN_19 = 3'h4 == _GEN_4 ? _source_WIRE_4 : _GEN_18; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire [2:0] _source_WIRE_5 = cams_5_io_key; // @[SourceA.scala 71:22 SourceA.scala 71:22]
  wire [2:0] _GEN_20 = 3'h5 == _GEN_4 ? _source_WIRE_5 : _GEN_19; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire [2:0] _source_WIRE_6 = cams_6_io_key; // @[SourceA.scala 71:22 SourceA.scala 71:22]
  wire [2:0] _GEN_21 = 3'h6 == _GEN_4 ? _source_WIRE_6 : _GEN_20; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire [2:0] _source_WIRE_7 = cams_7_io_key; // @[SourceA.scala 71:22 SourceA.scala 71:22]
  wire [2:0] _GEN_22 = 3'h7 == _GEN_4 ? _source_WIRE_7 : _GEN_21; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire [2:0] _GEN_23 = a_first ? _GEN_22 : source_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire [7:0] a_sel = 8'h1 << _GEN_4; // @[OneHot.scala 58:35]
  wire [63:0] _extract_io_i_bits_address_T = q_legal ? q_address : 64'h1000; // @[Parameters.scala 138:10]
  wire [51:0] extract_io_i_bits_address_hi = _extract_io_i_bits_address_T[63:12]; // @[Parameters.scala 138:47]
  wire [11:0] extract_io_i_bits_address_lo = q_address[11:0]; // @[Parameters.scala 139:14]
  wire [63:0] _extract_io_i_bits_address_T_1 = {extract_io_i_bits_address_hi,extract_io_i_bits_address_lo}; // @[Cat.scala 30:58]
  wire  extract_io_i_bits_mask_sizeOH_shiftAmount = _GEN_3[0]; // @[OneHot.scala 64:49]
  wire [1:0] _extract_io_i_bits_mask_sizeOH_T_1 = 2'h1 << extract_io_i_bits_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] extract_io_i_bits_mask_sizeOH = _extract_io_i_bits_mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _extract_io_i_bits_mask_T = _GEN_3 >= 4'h2; // @[Misc.scala 205:21]
  wire  extract_io_i_bits_mask_size = extract_io_i_bits_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  extract_io_i_bits_mask_bit = _GEN_6[1]; // @[Misc.scala 209:26]
  wire  extract_io_i_bits_mask_nbit = ~extract_io_i_bits_mask_bit; // @[Misc.scala 210:20]
  wire  extract_io_i_bits_mask_acc = _extract_io_i_bits_mask_T | extract_io_i_bits_mask_size &
    extract_io_i_bits_mask_nbit; // @[Misc.scala 214:29]
  wire  extract_io_i_bits_mask_acc_1 = _extract_io_i_bits_mask_T | extract_io_i_bits_mask_size &
    extract_io_i_bits_mask_bit; // @[Misc.scala 214:29]
  wire  extract_io_i_bits_mask_size_1 = extract_io_i_bits_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  extract_io_i_bits_mask_bit_1 = _GEN_6[0]; // @[Misc.scala 209:26]
  wire  extract_io_i_bits_mask_nbit_1 = ~extract_io_i_bits_mask_bit_1; // @[Misc.scala 210:20]
  wire  extract_io_i_bits_mask_eq_2 = extract_io_i_bits_mask_nbit & extract_io_i_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  extract_io_i_bits_mask_lo_lo = extract_io_i_bits_mask_acc | extract_io_i_bits_mask_size_1 &
    extract_io_i_bits_mask_eq_2; // @[Misc.scala 214:29]
  wire  extract_io_i_bits_mask_eq_3 = extract_io_i_bits_mask_nbit & extract_io_i_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  extract_io_i_bits_mask_lo_hi = extract_io_i_bits_mask_acc | extract_io_i_bits_mask_size_1 &
    extract_io_i_bits_mask_eq_3; // @[Misc.scala 214:29]
  wire  extract_io_i_bits_mask_eq_4 = extract_io_i_bits_mask_bit & extract_io_i_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  extract_io_i_bits_mask_hi_lo = extract_io_i_bits_mask_acc_1 | extract_io_i_bits_mask_size_1 &
    extract_io_i_bits_mask_eq_4; // @[Misc.scala 214:29]
  wire  extract_io_i_bits_mask_eq_5 = extract_io_i_bits_mask_bit & extract_io_i_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  extract_io_i_bits_mask_hi_hi = extract_io_i_bits_mask_acc_1 | extract_io_i_bits_mask_size_1 &
    extract_io_i_bits_mask_eq_5; // @[Misc.scala 214:29]
  wire [1:0] extract_io_i_bits_mask_lo = {extract_io_i_bits_mask_lo_hi,extract_io_i_bits_mask_lo_lo}; // @[Cat.scala 30:58]
  wire [1:0] extract_io_i_bits_mask_hi = {extract_io_i_bits_mask_hi_hi,extract_io_i_bits_mask_hi_lo}; // @[Cat.scala 30:58]
  wire  _source_ok_WIRE_0 = cams_0_io_alloc_ready; // @[SourceA.scala 70:22 SourceA.scala 70:22]
  wire  _source_ok_WIRE_1 = cams_1_io_alloc_ready; // @[SourceA.scala 70:22 SourceA.scala 70:22]
  wire  _GEN_25 = 3'h1 == _GEN_4 ? _source_ok_WIRE_1 : _source_ok_WIRE_0; // @[SourceA.scala 89:26 SourceA.scala 89:26]
  wire  _source_ok_WIRE_2 = cams_2_io_alloc_ready; // @[SourceA.scala 70:22 SourceA.scala 70:22]
  wire  _GEN_26 = 3'h2 == _GEN_4 ? _source_ok_WIRE_2 : _GEN_25; // @[SourceA.scala 89:26 SourceA.scala 89:26]
  wire  _source_ok_WIRE_3 = cams_3_io_alloc_ready; // @[SourceA.scala 70:22 SourceA.scala 70:22]
  wire  _GEN_27 = 3'h3 == _GEN_4 ? _source_ok_WIRE_3 : _GEN_26; // @[SourceA.scala 89:26 SourceA.scala 89:26]
  wire  _source_ok_WIRE_4 = cams_4_io_alloc_ready; // @[SourceA.scala 70:22 SourceA.scala 70:22]
  wire  _GEN_28 = 3'h4 == _GEN_4 ? _source_ok_WIRE_4 : _GEN_27; // @[SourceA.scala 89:26 SourceA.scala 89:26]
  wire  _source_ok_WIRE_5 = cams_5_io_alloc_ready; // @[SourceA.scala 70:22 SourceA.scala 70:22]
  wire  _GEN_29 = 3'h5 == _GEN_4 ? _source_ok_WIRE_5 : _GEN_28; // @[SourceA.scala 89:26 SourceA.scala 89:26]
  wire  _source_ok_WIRE_6 = cams_6_io_alloc_ready; // @[SourceA.scala 70:22 SourceA.scala 70:22]
  wire  _GEN_30 = 3'h6 == _GEN_4 ? _source_ok_WIRE_6 : _GEN_29; // @[SourceA.scala 89:26 SourceA.scala 89:26]
  wire  _source_ok_WIRE_7 = cams_7_io_alloc_ready; // @[SourceA.scala 70:22 SourceA.scala 70:22]
  wire  _GEN_31 = 3'h7 == _GEN_4 ? _source_ok_WIRE_7 : _GEN_30; // @[SourceA.scala 89:26 SourceA.scala 89:26]
  wire  stall = a_first & ~_GEN_31; // @[SourceA.scala 89:23]
  wire  xmit = q_last | state == 2'h3; // @[SourceA.scala 90:21]
  wire  _extract_io_i_valid_T = ~stall; // @[SourceA.scala 91:29]
  wire [2:0] d_clDomain = io_d_tlSource_bits[5:3]; // @[SourceA.scala 99:39]
  wire [7:0] d_sel = 8'h1 << d_clDomain; // @[OneHot.scala 58:35]
  wire [15:0] _io_d_clSource_WIRE_0 = cams_0_io_data; // @[SourceA.scala 101:23 SourceA.scala 101:23]
  wire [15:0] _io_d_clSource_WIRE_1 = cams_1_io_data; // @[SourceA.scala 101:23 SourceA.scala 101:23]
  wire [15:0] _GEN_33 = 3'h1 == d_clDomain ? _io_d_clSource_WIRE_1 : _io_d_clSource_WIRE_0; // @[SourceA.scala 101:17 SourceA.scala 101:17]
  wire [15:0] _io_d_clSource_WIRE_2 = cams_2_io_data; // @[SourceA.scala 101:23 SourceA.scala 101:23]
  wire [15:0] _GEN_34 = 3'h2 == d_clDomain ? _io_d_clSource_WIRE_2 : _GEN_33; // @[SourceA.scala 101:17 SourceA.scala 101:17]
  wire [15:0] _io_d_clSource_WIRE_3 = cams_3_io_data; // @[SourceA.scala 101:23 SourceA.scala 101:23]
  wire [15:0] _GEN_35 = 3'h3 == d_clDomain ? _io_d_clSource_WIRE_3 : _GEN_34; // @[SourceA.scala 101:17 SourceA.scala 101:17]
  wire [15:0] _io_d_clSource_WIRE_4 = cams_4_io_data; // @[SourceA.scala 101:23 SourceA.scala 101:23]
  wire [15:0] _GEN_36 = 3'h4 == d_clDomain ? _io_d_clSource_WIRE_4 : _GEN_35; // @[SourceA.scala 101:17 SourceA.scala 101:17]
  wire [15:0] _io_d_clSource_WIRE_5 = cams_5_io_data; // @[SourceA.scala 101:23 SourceA.scala 101:23]
  wire [15:0] _GEN_37 = 3'h5 == d_clDomain ? _io_d_clSource_WIRE_5 : _GEN_36; // @[SourceA.scala 101:17 SourceA.scala 101:17]
  wire [15:0] _io_d_clSource_WIRE_6 = cams_6_io_data; // @[SourceA.scala 101:23 SourceA.scala 101:23]
  wire [15:0] _GEN_38 = 3'h6 == d_clDomain ? _io_d_clSource_WIRE_6 : _GEN_37; // @[SourceA.scala 101:17 SourceA.scala 101:17]
  wire [15:0] _io_d_clSource_WIRE_7 = cams_7_io_data; // @[SourceA.scala 101:23 SourceA.scala 101:23]
  CAM cams_0 ( // @[SourceA.scala 21:11]
    .clock(cams_0_clock),
    .reset(cams_0_reset),
    .io_alloc_ready(cams_0_io_alloc_ready),
    .io_alloc_valid(cams_0_io_alloc_valid),
    .io_alloc_bits(cams_0_io_alloc_bits),
    .io_key(cams_0_io_key),
    .io_free_valid(cams_0_io_free_valid),
    .io_free_bits(cams_0_io_free_bits),
    .io_data(cams_0_io_data)
  );
  CAM cams_1 ( // @[SourceA.scala 21:11]
    .clock(cams_1_clock),
    .reset(cams_1_reset),
    .io_alloc_ready(cams_1_io_alloc_ready),
    .io_alloc_valid(cams_1_io_alloc_valid),
    .io_alloc_bits(cams_1_io_alloc_bits),
    .io_key(cams_1_io_key),
    .io_free_valid(cams_1_io_free_valid),
    .io_free_bits(cams_1_io_free_bits),
    .io_data(cams_1_io_data)
  );
  CAM cams_2 ( // @[SourceA.scala 21:11]
    .clock(cams_2_clock),
    .reset(cams_2_reset),
    .io_alloc_ready(cams_2_io_alloc_ready),
    .io_alloc_valid(cams_2_io_alloc_valid),
    .io_alloc_bits(cams_2_io_alloc_bits),
    .io_key(cams_2_io_key),
    .io_free_valid(cams_2_io_free_valid),
    .io_free_bits(cams_2_io_free_bits),
    .io_data(cams_2_io_data)
  );
  CAM cams_3 ( // @[SourceA.scala 21:11]
    .clock(cams_3_clock),
    .reset(cams_3_reset),
    .io_alloc_ready(cams_3_io_alloc_ready),
    .io_alloc_valid(cams_3_io_alloc_valid),
    .io_alloc_bits(cams_3_io_alloc_bits),
    .io_key(cams_3_io_key),
    .io_free_valid(cams_3_io_free_valid),
    .io_free_bits(cams_3_io_free_bits),
    .io_data(cams_3_io_data)
  );
  CAM cams_4 ( // @[SourceA.scala 21:11]
    .clock(cams_4_clock),
    .reset(cams_4_reset),
    .io_alloc_ready(cams_4_io_alloc_ready),
    .io_alloc_valid(cams_4_io_alloc_valid),
    .io_alloc_bits(cams_4_io_alloc_bits),
    .io_key(cams_4_io_key),
    .io_free_valid(cams_4_io_free_valid),
    .io_free_bits(cams_4_io_free_bits),
    .io_data(cams_4_io_data)
  );
  CAM cams_5 ( // @[SourceA.scala 21:11]
    .clock(cams_5_clock),
    .reset(cams_5_reset),
    .io_alloc_ready(cams_5_io_alloc_ready),
    .io_alloc_valid(cams_5_io_alloc_valid),
    .io_alloc_bits(cams_5_io_alloc_bits),
    .io_key(cams_5_io_key),
    .io_free_valid(cams_5_io_free_valid),
    .io_free_bits(cams_5_io_free_bits),
    .io_data(cams_5_io_data)
  );
  CAM cams_6 ( // @[SourceA.scala 21:11]
    .clock(cams_6_clock),
    .reset(cams_6_reset),
    .io_alloc_ready(cams_6_io_alloc_ready),
    .io_alloc_valid(cams_6_io_alloc_valid),
    .io_alloc_bits(cams_6_io_alloc_bits),
    .io_key(cams_6_io_key),
    .io_free_valid(cams_6_io_free_valid),
    .io_free_bits(cams_6_io_free_bits),
    .io_data(cams_6_io_data)
  );
  CAM cams_7 ( // @[SourceA.scala 21:11]
    .clock(cams_7_clock),
    .reset(cams_7_reset),
    .io_alloc_ready(cams_7_io_alloc_ready),
    .io_alloc_valid(cams_7_io_alloc_valid),
    .io_alloc_bits(cams_7_io_alloc_bits),
    .io_key(cams_7_io_key),
    .io_free_valid(cams_7_io_free_valid),
    .io_free_bits(cams_7_io_free_bits),
    .io_data(cams_7_io_data)
  );
  ParitalExtractor extract ( // @[SourceA.scala 75:23]
    .clock(extract_clock),
    .reset(extract_reset),
    .io_last(extract_io_last),
    .io_i_ready(extract_io_i_ready),
    .io_i_valid(extract_io_i_valid),
    .io_i_bits_opcode(extract_io_i_bits_opcode),
    .io_i_bits_param(extract_io_i_bits_param),
    .io_i_bits_size(extract_io_i_bits_size),
    .io_i_bits_source(extract_io_i_bits_source),
    .io_i_bits_address(extract_io_i_bits_address),
    .io_i_bits_mask(extract_io_i_bits_mask),
    .io_i_bits_data(extract_io_i_bits_data),
    .io_o_ready(extract_io_o_ready),
    .io_o_valid(extract_io_o_valid),
    .io_o_bits_opcode(extract_io_o_bits_opcode),
    .io_o_bits_param(extract_io_o_bits_param),
    .io_o_bits_size(extract_io_o_bits_size),
    .io_o_bits_source(extract_io_o_bits_source),
    .io_o_bits_address(extract_io_o_bits_address),
    .io_o_bits_mask(extract_io_o_bits_mask),
    .io_o_bits_data(extract_io_o_bits_data)
  );
  assign io_a_valid = extract_io_o_valid; // @[SourceA.scala 76:8]
  assign io_a_bits_opcode = extract_io_o_bits_opcode; // @[SourceA.scala 76:8]
  assign io_a_bits_param = extract_io_o_bits_param; // @[SourceA.scala 76:8]
  assign io_a_bits_size = extract_io_o_bits_size; // @[SourceA.scala 76:8]
  assign io_a_bits_source = extract_io_o_bits_source; // @[SourceA.scala 76:8]
  assign io_a_bits_address = extract_io_o_bits_address; // @[SourceA.scala 76:8]
  assign io_a_bits_mask = extract_io_o_bits_mask; // @[SourceA.scala 76:8]
  assign io_a_bits_data = extract_io_o_bits_data; // @[SourceA.scala 76:8]
  assign io_q_ready = extract_io_i_ready & _extract_io_i_valid_T | ~xmit; // @[SourceA.scala 92:37]
  assign io_d_clSource = 3'h7 == d_clDomain ? _io_d_clSource_WIRE_7 : _GEN_38; // @[SourceA.scala 101:17 SourceA.scala 101:17]
  assign cams_0_clock = clock;
  assign cams_0_reset = reset;
  assign cams_0_io_alloc_valid = a_sel[0] & a_first & xmit & io_q_valid & extract_io_i_ready; // @[SourceA.scala 94:64]
  assign cams_0_io_alloc_bits = enable ? source : r_5; // @[SourceA.scala 33:8]
  assign cams_0_io_free_valid = io_d_tlSource_valid & d_sel[0]; // @[SourceA.scala 104:46]
  assign cams_0_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceA.scala 103:23]
  assign cams_1_clock = clock;
  assign cams_1_reset = reset;
  assign cams_1_io_alloc_valid = a_sel[1] & a_first & xmit & io_q_valid & extract_io_i_ready; // @[SourceA.scala 94:64]
  assign cams_1_io_alloc_bits = enable ? source : r_5; // @[SourceA.scala 33:8]
  assign cams_1_io_free_valid = io_d_tlSource_valid & d_sel[1]; // @[SourceA.scala 104:46]
  assign cams_1_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceA.scala 103:23]
  assign cams_2_clock = clock;
  assign cams_2_reset = reset;
  assign cams_2_io_alloc_valid = a_sel[2] & a_first & xmit & io_q_valid & extract_io_i_ready; // @[SourceA.scala 94:64]
  assign cams_2_io_alloc_bits = enable ? source : r_5; // @[SourceA.scala 33:8]
  assign cams_2_io_free_valid = io_d_tlSource_valid & d_sel[2]; // @[SourceA.scala 104:46]
  assign cams_2_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceA.scala 103:23]
  assign cams_3_clock = clock;
  assign cams_3_reset = reset;
  assign cams_3_io_alloc_valid = a_sel[3] & a_first & xmit & io_q_valid & extract_io_i_ready; // @[SourceA.scala 94:64]
  assign cams_3_io_alloc_bits = enable ? source : r_5; // @[SourceA.scala 33:8]
  assign cams_3_io_free_valid = io_d_tlSource_valid & d_sel[3]; // @[SourceA.scala 104:46]
  assign cams_3_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceA.scala 103:23]
  assign cams_4_clock = clock;
  assign cams_4_reset = reset;
  assign cams_4_io_alloc_valid = a_sel[4] & a_first & xmit & io_q_valid & extract_io_i_ready; // @[SourceA.scala 94:64]
  assign cams_4_io_alloc_bits = enable ? source : r_5; // @[SourceA.scala 33:8]
  assign cams_4_io_free_valid = io_d_tlSource_valid & d_sel[4]; // @[SourceA.scala 104:46]
  assign cams_4_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceA.scala 103:23]
  assign cams_5_clock = clock;
  assign cams_5_reset = reset;
  assign cams_5_io_alloc_valid = a_sel[5] & a_first & xmit & io_q_valid & extract_io_i_ready; // @[SourceA.scala 94:64]
  assign cams_5_io_alloc_bits = enable ? source : r_5; // @[SourceA.scala 33:8]
  assign cams_5_io_free_valid = io_d_tlSource_valid & d_sel[5]; // @[SourceA.scala 104:46]
  assign cams_5_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceA.scala 103:23]
  assign cams_6_clock = clock;
  assign cams_6_reset = reset;
  assign cams_6_io_alloc_valid = a_sel[6] & a_first & xmit & io_q_valid & extract_io_i_ready; // @[SourceA.scala 94:64]
  assign cams_6_io_alloc_bits = enable ? source : r_5; // @[SourceA.scala 33:8]
  assign cams_6_io_free_valid = io_d_tlSource_valid & d_sel[6]; // @[SourceA.scala 104:46]
  assign cams_6_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceA.scala 103:23]
  assign cams_7_clock = clock;
  assign cams_7_reset = reset;
  assign cams_7_io_alloc_valid = a_sel[7] & a_first & xmit & io_q_valid & extract_io_i_ready; // @[SourceA.scala 94:64]
  assign cams_7_io_alloc_bits = enable ? source : r_5; // @[SourceA.scala 33:8]
  assign cams_7_io_free_valid = io_d_tlSource_valid & d_sel[7]; // @[SourceA.scala 104:46]
  assign cams_7_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceA.scala 103:23]
  assign extract_clock = clock;
  assign extract_reset = reset;
  assign extract_io_last = q_last_count == 5'h1 | q_last_first & q_last_beats_a == 5'h0; // @[Parameters.scala 129:35]
  assign extract_io_i_valid = io_q_valid & ~stall & xmit; // @[SourceA.scala 91:37]
  assign extract_io_i_bits_opcode = enable ? opcode : r_1; // @[SourceA.scala 33:8]
  assign extract_io_i_bits_param = enable ? param : r_2; // @[SourceA.scala 33:8]
  assign extract_io_i_bits_size = _GEN_3[2:0]; // @[SourceA.scala 82:18]
  assign extract_io_i_bits_source = {_GEN_4,_GEN_23}; // @[Cat.scala 30:58]
  assign extract_io_i_bits_address = _extract_io_i_bits_address_T_1[31:0]; // @[SourceA.scala 84:18]
  assign extract_io_i_bits_mask = {extract_io_i_bits_mask_hi,extract_io_i_bits_mask_lo}; // @[Cat.scala 30:58]
  assign extract_io_i_bits_data = io_q_bits; // @[SourceA.scala 86:18]
  assign extract_io_o_ready = io_a_ready; // @[SourceA.scala 76:8]
  always @(posedge clock) begin
    if (reset) begin // @[SourceA.scala 25:22]
      state <= 2'h0; // @[SourceA.scala 25:22]
    end else if (_q_last_T) begin // @[SourceA.scala 48:22]
      if (_T_2) begin // @[Conditional.scala 40:58]
        state <= 2'h1; // @[SourceA.scala 50:31]
      end else if (_T_3) begin // @[Conditional.scala 39:67]
        state <= 2'h2; // @[SourceA.scala 51:31]
      end else begin
        state <= _GEN_11;
      end
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_1 <= opcode; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_2 <= param; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_3 <= size; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_4 <= domain; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_5 <= source; // @[Reg.scala 16:23]
    end
    if (q_address0_enable) begin // @[Reg.scala 16:19]
      q_address0_r <= io_q_bits; // @[Reg.scala 16:23]
    end
    if (q_address1_enable) begin // @[Reg.scala 16:19]
      q_address1_r <= io_q_bits; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Parameters.scala 126:24]
      q_last_count <= 5'h0; // @[Parameters.scala 126:24]
    end else if (_q_last_T) begin // @[Parameters.scala 130:21]
      if (q_last_first) begin // @[Parameters.scala 130:35]
        q_last_count <= q_last_beats_a;
      end else begin
        q_last_count <= _q_last_count_T_1;
      end
    end
    if (_q_last_T) begin // @[Reg.scala 16:19]
      a_first <= _a_first_T; // @[Reg.scala 16:23]
    end
    if (a_first) begin // @[Reg.scala 16:19]
      if (3'h7 == _GEN_4) begin // @[Reg.scala 16:23]
        source_r <= _source_WIRE_7; // @[Reg.scala 16:23]
      end else if (3'h6 == _GEN_4) begin // @[Reg.scala 16:23]
        source_r <= _source_WIRE_6; // @[Reg.scala 16:23]
      end else if (3'h5 == _GEN_4) begin // @[Reg.scala 16:23]
        source_r <= _source_WIRE_5; // @[Reg.scala 16:23]
      end else begin
        source_r <= _GEN_19;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  r_4 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  r_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  q_address0_r = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  q_address1_r = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  q_last_count = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  a_first = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  source_r = _RAND_10[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ParitalExtractor_1(
  input        clock,
  input        reset,
  input        io_last,
  output       io_i_ready,
  input        io_i_valid,
  input  [2:0] io_i_bits_opcode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] state; // @[Partial.scala 29:23]
  wire  enable = io_i_bits_opcode == 3'h1; // @[Partial.scala 31:25]
  wire  empty = state == 4'h0; // @[Partial.scala 32:22]
  wire  _T = io_i_ready & io_i_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _state_T_1 = state - 4'h1; // @[Partial.scala 48:22]
  wire [3:0] _GEN_2 = empty ? 4'h8 : _state_T_1; // @[Partial.scala 49:22 Partial.scala 49:30 Partial.scala 48:13]
  assign io_i_ready = enable & empty; // @[Partial.scala 34:17 Partial.scala 17:8]
  always @(posedge clock) begin
    if (reset) begin // @[Partial.scala 29:23]
      state <= 4'h0; // @[Partial.scala 29:23]
    end else if (enable) begin // @[Partial.scala 34:17]
      if (_T) begin // @[Partial.scala 46:24]
        if (io_last) begin // @[Partial.scala 50:22]
          state <= 4'h0; // @[Partial.scala 50:30]
        end else begin
          state <= _GEN_2;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SourceB(
  input         clock,
  input         reset,
  output        io_q_ready,
  input         io_q_valid,
  input  [31:0] io_q_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  extract_clock; // @[SourceB.scala 53:23]
  wire  extract_reset; // @[SourceB.scala 53:23]
  wire  extract_io_last; // @[SourceB.scala 53:23]
  wire  extract_io_i_ready; // @[SourceB.scala 53:23]
  wire  extract_io_i_valid; // @[SourceB.scala 53:23]
  wire [2:0] extract_io_i_bits_opcode; // @[SourceB.scala 53:23]
  reg [1:0] state; // @[SourceB.scala 20:22]
  wire [2:0] opcode = io_q_bits[5:3]; // @[Parameters.scala 92:19]
  wire [3:0] size = io_q_bits[12:9]; // @[Parameters.scala 94:19]
  wire  enable = state == 2'h0; // @[SourceB.scala 27:24]
  reg [2:0] r_1; // @[Reg.scala 15:16]
  wire [2:0] _GEN_1 = enable ? opcode : r_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [4:0] q_last_count; // @[Parameters.scala 126:24]
  wire [2:0] q_last_beats_beats_shiftAmount = size[2:0]; // @[OneHot.scala 64:49]
  wire [7:0] _q_last_beats_beats_T_1 = 8'h1 << q_last_beats_beats_shiftAmount; // @[OneHot.scala 65:12]
  wire [3:0] q_last_beats_beats_hi = _q_last_beats_beats_T_1[6:3]; // @[Parameters.scala 102:62]
  wire  q_last_beats_beats_lo = size <= 4'h2; // @[Parameters.scala 102:83]
  wire [4:0] q_last_beats_beats = {q_last_beats_beats_hi,q_last_beats_beats_lo}; // @[Cat.scala 30:58]
  wire  q_last_beats_masks_hi = _q_last_beats_beats_T_1[6]; // @[Parameters.scala 107:62]
  wire  q_last_beats_masks_lo = size <= 4'h5; // @[Parameters.scala 107:83]
  wire [1:0] q_last_beats_masks = {q_last_beats_masks_hi,q_last_beats_masks_lo}; // @[Cat.scala 30:58]
  wire  q_last_beats_partial = opcode == 3'h1; // @[Parameters.scala 115:26]
  wire [4:0] _q_last_beats_a_T_1 = opcode[2] ? 5'h0 : q_last_beats_beats; // @[Parameters.scala 116:16]
  wire [4:0] _q_last_beats_a_T_3 = _q_last_beats_a_T_1 + 5'h2; // @[Parameters.scala 116:44]
  wire [1:0] _q_last_beats_a_T_4 = q_last_beats_partial ? q_last_beats_masks : 2'h0; // @[Parameters.scala 116:59]
  wire [4:0] _GEN_15 = {{3'd0}, _q_last_beats_a_T_4}; // @[Parameters.scala 116:54]
  wire [4:0] q_last_beats_a = _q_last_beats_a_T_3 + _GEN_15; // @[Parameters.scala 116:54]
  wire  q_last_first = q_last_count == 5'h0; // @[Parameters.scala 128:23]
  wire  q_last = q_last_count == 5'h1 | q_last_first & q_last_beats_a == 5'h0; // @[Parameters.scala 129:35]
  wire  _q_last_T = io_q_ready & io_q_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _q_last_count_T_1 = q_last_count - 5'h1; // @[Parameters.scala 130:56]
  wire  q_hasData = ~_GEN_1[2]; // @[SourceB.scala 40:19]
  wire  _T_4 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T = q_hasData ? 2'h3 : 2'h0; // @[SourceB.scala 47:37]
  wire  _T_7 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T_2 = ~q_last ? 2'h3 : 2'h0; // @[SourceB.scala 48:37]
  wire [1:0] _GEN_10 = _T_7 ? _state_T_2 : state; // @[Conditional.scala 39:67 SourceB.scala 48:31 SourceB.scala 20:22]
  wire [1:0] _GEN_11 = _T_6 ? _state_T : _GEN_10; // @[Conditional.scala 39:67 SourceB.scala 47:31]
  wire  xmit = q_last | state == 2'h3; // @[SourceB.scala 67:21]
  ParitalExtractor_1 extract ( // @[SourceB.scala 53:23]
    .clock(extract_clock),
    .reset(extract_reset),
    .io_last(extract_io_last),
    .io_i_ready(extract_io_i_ready),
    .io_i_valid(extract_io_i_valid),
    .io_i_bits_opcode(extract_io_i_bits_opcode)
  );
  assign io_q_ready = extract_io_i_ready | ~xmit; // @[SourceB.scala 69:25]
  assign extract_clock = clock;
  assign extract_reset = reset;
  assign extract_io_last = q_last_count == 5'h1 | q_last_first & q_last_beats_a == 5'h0; // @[Parameters.scala 129:35]
  assign extract_io_i_valid = io_q_valid & xmit; // @[SourceB.scala 68:25]
  assign extract_io_i_bits_opcode = enable ? opcode : r_1; // @[SourceB.scala 28:8]
  always @(posedge clock) begin
    if (reset) begin // @[SourceB.scala 20:22]
      state <= 2'h0; // @[SourceB.scala 20:22]
    end else if (_q_last_T) begin // @[SourceB.scala 43:22]
      if (_T_4) begin // @[Conditional.scala 40:58]
        state <= 2'h1; // @[SourceB.scala 45:31]
      end else if (_T_5) begin // @[Conditional.scala 39:67]
        state <= 2'h2; // @[SourceB.scala 46:31]
      end else begin
        state <= _GEN_11;
      end
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_1 <= opcode; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Parameters.scala 126:24]
      q_last_count <= 5'h0; // @[Parameters.scala 126:24]
    end else if (_q_last_T) begin // @[Parameters.scala 130:21]
      if (q_last_first) begin // @[Parameters.scala 130:35]
        q_last_count <= q_last_beats_a;
      end else begin
        q_last_count <= _q_last_count_T_1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  q_last_count = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CAM_8(
  input         clock,
  input         reset,
  output        io_alloc_ready,
  input         io_alloc_valid,
  input  [15:0] io_alloc_bits,
  output [2:0]  io_key,
  input         io_free_valid,
  input  [2:0]  io_free_bits,
  output [15:0] io_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] data [0:7]; // @[CAM.scala 22:17]
  wire [15:0] data_io_data_MPORT_data; // @[CAM.scala 22:17]
  wire [2:0] data_io_data_MPORT_addr; // @[CAM.scala 22:17]
  wire [15:0] data_MPORT_data; // @[CAM.scala 22:17]
  wire [2:0] data_MPORT_addr; // @[CAM.scala 22:17]
  wire  data_MPORT_mask; // @[CAM.scala 22:17]
  wire  data_MPORT_en; // @[CAM.scala 22:17]
  reg [7:0] free; // @[CAM.scala 21:21]
  wire [8:0] _free_sel_T = {free, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _free_sel_T_2 = free | _free_sel_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _free_sel_T_3 = {_free_sel_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _free_sel_T_5 = _free_sel_T_2 | _free_sel_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _free_sel_T_6 = {_free_sel_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _free_sel_T_8 = _free_sel_T_5 | _free_sel_T_6[7:0]; // @[package.scala 244:43]
  wire [8:0] _free_sel_T_10 = {_free_sel_T_8, 1'h0}; // @[CAM.scala 24:39]
  wire [8:0] _free_sel_T_11 = ~_free_sel_T_10; // @[CAM.scala 24:18]
  wire [8:0] _GEN_5 = {{1'd0}, free}; // @[CAM.scala 24:45]
  wire [8:0] free_sel = _free_sel_T_11 & _GEN_5; // @[CAM.scala 24:45]
  wire [3:0] io_key_hi = free_sel[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] io_key_lo = free_sel[3:0]; // @[OneHot.scala 31:18]
  wire  io_key_hi_1 = |io_key_hi; // @[OneHot.scala 32:14]
  wire [3:0] _io_key_T = io_key_hi | io_key_lo; // @[OneHot.scala 32:28]
  wire [1:0] io_key_hi_2 = _io_key_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_key_lo_1 = _io_key_T[1:0]; // @[OneHot.scala 31:18]
  wire  io_key_hi_3 = |io_key_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _io_key_T_1 = io_key_hi_2 | io_key_lo_1; // @[OneHot.scala 32:28]
  wire  io_key_lo_2 = _io_key_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] io_key_lo_3 = {io_key_hi_3,io_key_lo_2}; // @[Cat.scala 30:58]
  wire  _T = io_alloc_ready & io_alloc_valid; // @[Decoupled.scala 40:37]
  wire  bypass = _T & io_free_bits == io_key; // @[CAM.scala 31:32]
  wire [8:0] clr = _T ? free_sel : 9'h0; // @[CAM.scala 35:16]
  wire [7:0] _set_T = 8'h1 << io_free_bits; // @[OneHot.scala 58:35]
  wire [7:0] set = io_free_valid ? _set_T : 8'h0; // @[CAM.scala 36:16]
  wire [8:0] _free_T = ~clr; // @[CAM.scala 37:19]
  wire [8:0] _free_T_1 = _GEN_5 & _free_T; // @[CAM.scala 37:17]
  wire [8:0] _GEN_7 = {{1'd0}, set}; // @[CAM.scala 37:25]
  wire [8:0] _free_T_2 = _free_T_1 | _GEN_7; // @[CAM.scala 37:25]
  assign data_io_data_MPORT_addr = io_free_bits;
  assign data_io_data_MPORT_data = data[data_io_data_MPORT_addr]; // @[CAM.scala 22:17]
  assign data_MPORT_data = io_alloc_bits;
  assign data_MPORT_addr = io_key;
  assign data_MPORT_mask = 1'h1;
  assign data_MPORT_en = io_alloc_ready & io_alloc_valid;
  assign io_alloc_ready = |free; // @[CAM.scala 27:26]
  assign io_key = {io_key_hi_1,io_key_lo_3}; // @[Cat.scala 30:58]
  assign io_data = bypass ? io_alloc_bits : data_io_data_MPORT_data; // @[CAM.scala 32:17]
  always @(posedge clock) begin
    if(data_MPORT_en & data_MPORT_mask) begin
      data[data_MPORT_addr] <= data_MPORT_data; // @[CAM.scala 22:17]
    end
    if (reset) begin // @[CAM.scala 21:21]
      free <= 8'hff; // @[CAM.scala 21:21]
    end else begin
      free <= _free_T_2[7:0]; // @[CAM.scala 37:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  free = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SourceC(
  input         clock,
  input         reset,
  input         io_c_ready,
  output        io_c_valid,
  output [2:0]  io_c_bits_opcode,
  output [2:0]  io_c_bits_param,
  output [2:0]  io_c_bits_size,
  output [5:0]  io_c_bits_source,
  output [31:0] io_c_bits_address,
  output        io_q_ready,
  input         io_q_valid,
  input  [31:0] io_q_bits,
  input         io_d_tlSource_valid,
  input  [5:0]  io_d_tlSource_bits,
  output [15:0] io_d_clSource
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  cam_clock; // @[SourceC.scala 20:19]
  wire  cam_reset; // @[SourceC.scala 20:19]
  wire  cam_io_alloc_ready; // @[SourceC.scala 20:19]
  wire  cam_io_alloc_valid; // @[SourceC.scala 20:19]
  wire [15:0] cam_io_alloc_bits; // @[SourceC.scala 20:19]
  wire [2:0] cam_io_key; // @[SourceC.scala 20:19]
  wire  cam_io_free_valid; // @[SourceC.scala 20:19]
  wire [2:0] cam_io_free_bits; // @[SourceC.scala 20:19]
  wire [15:0] cam_io_data; // @[SourceC.scala 20:19]
  reg [1:0] state; // @[SourceC.scala 23:22]
  wire [2:0] opcode = io_q_bits[5:3]; // @[Parameters.scala 92:19]
  wire [2:0] param = io_q_bits[8:6]; // @[Parameters.scala 93:19]
  wire [3:0] size = io_q_bits[12:9]; // @[Parameters.scala 94:19]
  wire [15:0] source = io_q_bits[31:16]; // @[Parameters.scala 96:19]
  wire  enable = state == 2'h0; // @[SourceC.scala 30:24]
  reg [2:0] r_1; // @[Reg.scala 15:16]
  wire [2:0] _GEN_1 = enable ? opcode : r_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [2:0] r_2; // @[Reg.scala 15:16]
  reg [3:0] r_3; // @[Reg.scala 15:16]
  wire [3:0] _GEN_3 = enable ? size : r_3; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [15:0] r_5; // @[Reg.scala 15:16]
  wire  q_address0_enable = state == 2'h1; // @[SourceC.scala 30:24]
  reg [31:0] q_address0_r; // @[Reg.scala 15:16]
  wire [31:0] _GEN_6 = q_address0_enable ? io_q_bits : q_address0_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire  q_address1_enable = state == 2'h2; // @[SourceC.scala 30:24]
  reg [31:0] q_address1_r; // @[Reg.scala 15:16]
  wire [31:0] _GEN_7 = q_address1_enable ? io_q_bits : q_address1_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [4:0] q_last_count; // @[Parameters.scala 126:24]
  wire [2:0] q_last_beats_beats_shiftAmount = size[2:0]; // @[OneHot.scala 64:49]
  wire [7:0] _q_last_beats_beats_T_1 = 8'h1 << q_last_beats_beats_shiftAmount; // @[OneHot.scala 65:12]
  wire [3:0] q_last_beats_beats_hi = _q_last_beats_beats_T_1[6:3]; // @[Parameters.scala 102:62]
  wire  q_last_beats_beats_lo = size <= 4'h2; // @[Parameters.scala 102:83]
  wire [4:0] q_last_beats_beats = {q_last_beats_beats_hi,q_last_beats_beats_lo}; // @[Cat.scala 30:58]
  wire [4:0] _q_last_beats_c_T_1 = opcode[0] ? q_last_beats_beats : 5'h0; // @[Parameters.scala 118:16]
  wire [4:0] q_last_beats_c = _q_last_beats_c_T_1 + 5'h2; // @[Parameters.scala 118:44]
  wire  q_last_first = q_last_count == 5'h0; // @[Parameters.scala 128:23]
  wire  q_last = q_last_count == 5'h1 | q_last_first & q_last_beats_c == 5'h0; // @[Parameters.scala 129:35]
  wire  _q_last_T = io_q_ready & io_q_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _q_last_count_T_1 = q_last_count - 5'h1; // @[Parameters.scala 130:56]
  wire  q_hasData = _GEN_1[0]; // @[SourceC.scala 43:27]
  wire  _c_first_T = state != 2'h3; // @[SourceC.scala 44:33]
  reg  c_first; // @[Reg.scala 15:16]
  wire  _T_3 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T = q_hasData ? 2'h3 : 2'h0; // @[SourceC.scala 50:37]
  wire  _T_6 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _state_T_2 = ~q_last ? 2'h3 : 2'h0; // @[SourceC.scala 51:37]
  wire [1:0] _GEN_10 = _T_6 ? _state_T_2 : state; // @[Conditional.scala 39:67 SourceC.scala 51:31 SourceC.scala 23:22]
  wire [1:0] _GEN_11 = _T_5 ? _state_T : _GEN_10; // @[Conditional.scala 39:67 SourceC.scala 50:31]
  wire [63:0] q_address = {_GEN_7,_GEN_6}; // @[Cat.scala 30:58]
  wire [63:0] _exists_T = q_address ^ 64'h10000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_1 = {1'b0,$signed(_exists_T)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_3 = $signed(_exists_T_1) & -65'sh10000000; // @[Parameters.scala 137:52]
  wire  _exists_T_4 = $signed(_exists_T_3) == 65'sh0; // @[Parameters.scala 137:67]
  wire [63:0] _exists_T_5 = q_address ^ 64'h20000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_6 = {1'b0,$signed(_exists_T_5)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_8 = $signed(_exists_T_6) & -65'sh20000000; // @[Parameters.scala 137:52]
  wire  _exists_T_9 = $signed(_exists_T_8) == 65'sh0; // @[Parameters.scala 137:67]
  wire [63:0] _exists_T_10 = q_address ^ 64'h40000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_11 = {1'b0,$signed(_exists_T_10)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_13 = $signed(_exists_T_11) & -65'sh40000000; // @[Parameters.scala 137:52]
  wire  _exists_T_14 = $signed(_exists_T_13) == 65'sh0; // @[Parameters.scala 137:67]
  wire [63:0] _exists_T_15 = q_address ^ 64'h80000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_16 = {1'b0,$signed(_exists_T_15)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_18 = $signed(_exists_T_16) & -65'sh40000000; // @[Parameters.scala 137:52]
  wire  _exists_T_19 = $signed(_exists_T_18) == 65'sh0; // @[Parameters.scala 137:67]
  wire [63:0] _exists_T_20 = q_address ^ 64'hc0000000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_21 = {1'b0,$signed(_exists_T_20)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_23 = $signed(_exists_T_21) & -65'sh20000000; // @[Parameters.scala 137:52]
  wire  _exists_T_24 = $signed(_exists_T_23) == 65'sh0; // @[Parameters.scala 137:67]
  wire  _exists_T_28 = _exists_T_4 | _exists_T_9 | _exists_T_14 | _exists_T_19 | _exists_T_24; // @[Parameters.scala 598:92]
  wire [63:0] _exists_T_29 = q_address ^ 64'h1000; // @[Parameters.scala 137:31]
  wire [64:0] _exists_T_30 = {1'b0,$signed(_exists_T_29)}; // @[Parameters.scala 137:49]
  wire [64:0] _exists_T_32 = $signed(_exists_T_30) & -65'sh1000; // @[Parameters.scala 137:52]
  wire  _exists_T_33 = $signed(_exists_T_32) == 65'sh0; // @[Parameters.scala 137:67]
  wire  exists = _exists_T_28 | _exists_T_33; // @[Parameters.scala 622:64]
  wire [64:0] _writeOk_T_1 = {1'b0,$signed(q_address)}; // @[Parameters.scala 137:49]
  wire [64:0] _acquireOk_T_32 = $signed(_writeOk_T_1) & 65'shf0000000; // @[Parameters.scala 137:52]
  wire  acquireOk = $signed(_acquireOk_T_32) == 65'sh0; // @[Parameters.scala 137:67]
  wire  q_legal = exists & acquireOk; // @[SourceC.scala 63:51]
  wire  q_release = _GEN_1 == 3'h6 | _GEN_1 == 3'h7; // @[SourceC.scala 66:51]
  wire  source_ok = ~q_release | cam_io_alloc_ready; // @[SourceC.scala 67:30]
  reg [2:0] source_r; // @[Reg.scala 15:16]
  wire [2:0] _GEN_15 = c_first ? cam_io_key : source_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire [2:0] _io_c_bits_source_T = q_release ? _GEN_15 : 3'h0; // @[SourceC.scala 73:27]
  wire [63:0] _io_c_bits_address_T = q_legal ? q_address : 64'h1000; // @[Parameters.scala 138:10]
  wire [51:0] io_c_bits_address_hi = _io_c_bits_address_T[63:12]; // @[Parameters.scala 138:47]
  wire [11:0] io_c_bits_address_lo = q_address[11:0]; // @[Parameters.scala 139:14]
  wire [63:0] _io_c_bits_address_T_1 = {io_c_bits_address_hi,io_c_bits_address_lo}; // @[Cat.scala 30:58]
  wire  stall = c_first & ~source_ok; // @[SourceC.scala 78:23]
  wire  xmit = q_last | state == 2'h3; // @[SourceC.scala 79:21]
  wire  _io_c_valid_T = ~stall; // @[SourceC.scala 80:32]
  CAM_8 cam ( // @[SourceC.scala 20:19]
    .clock(cam_clock),
    .reset(cam_reset),
    .io_alloc_ready(cam_io_alloc_ready),
    .io_alloc_valid(cam_io_alloc_valid),
    .io_alloc_bits(cam_io_alloc_bits),
    .io_key(cam_io_key),
    .io_free_valid(cam_io_free_valid),
    .io_free_bits(cam_io_free_bits),
    .io_data(cam_io_data)
  );
  assign io_c_valid = io_q_valid & ~stall & xmit; // @[SourceC.scala 80:40]
  assign io_c_bits_opcode = enable ? opcode : r_1; // @[SourceC.scala 31:8]
  assign io_c_bits_param = enable ? param : r_2; // @[SourceC.scala 31:8]
  assign io_c_bits_size = _GEN_3[2:0]; // @[SourceC.scala 72:21]
  assign io_c_bits_source = {{3'd0}, _io_c_bits_source_T}; // @[SourceC.scala 73:27]
  assign io_c_bits_address = _io_c_bits_address_T_1[31:0]; // @[SourceC.scala 74:21]
  assign io_q_ready = io_c_ready & _io_c_valid_T | ~xmit; // @[SourceC.scala 81:40]
  assign io_d_clSource = cam_io_data; // @[SourceC.scala 86:17]
  assign cam_clock = clock;
  assign cam_reset = reset;
  assign cam_io_alloc_valid = q_release & c_first & xmit & io_q_valid & io_c_ready; // @[SourceC.scala 82:68]
  assign cam_io_alloc_bits = enable ? source : r_5; // @[SourceC.scala 31:8]
  assign cam_io_free_valid = io_d_tlSource_valid; // @[SourceC.scala 87:15]
  assign cam_io_free_bits = io_d_tlSource_bits[2:0]; // @[SourceC.scala 87:15]
  always @(posedge clock) begin
    if (reset) begin // @[SourceC.scala 23:22]
      state <= 2'h0; // @[SourceC.scala 23:22]
    end else if (_q_last_T) begin // @[SourceC.scala 46:22]
      if (_T_3) begin // @[Conditional.scala 40:58]
        state <= 2'h1; // @[SourceC.scala 48:31]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        state <= 2'h2; // @[SourceC.scala 49:31]
      end else begin
        state <= _GEN_11;
      end
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_1 <= opcode; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_2 <= param; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_3 <= size; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_5 <= source; // @[Reg.scala 16:23]
    end
    if (q_address0_enable) begin // @[Reg.scala 16:19]
      q_address0_r <= io_q_bits; // @[Reg.scala 16:23]
    end
    if (q_address1_enable) begin // @[Reg.scala 16:19]
      q_address1_r <= io_q_bits; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Parameters.scala 126:24]
      q_last_count <= 5'h0; // @[Parameters.scala 126:24]
    end else if (_q_last_T) begin // @[Parameters.scala 130:21]
      if (q_last_first) begin // @[Parameters.scala 130:35]
        q_last_count <= q_last_beats_c;
      end else begin
        q_last_count <= _q_last_count_T_1;
      end
    end
    if (_q_last_T) begin // @[Reg.scala 16:19]
      c_first <= _c_first_T; // @[Reg.scala 16:23]
    end
    if (c_first) begin // @[Reg.scala 16:19]
      source_r <= cam_io_key; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  r_5 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  q_address0_r = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  q_address1_r = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  q_last_count = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  c_first = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  source_r = _RAND_9[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CAM_9(
  input         clock,
  input         reset,
  output        io_alloc_ready,
  input         io_alloc_valid,
  input  [15:0] io_alloc_bits,
  output [4:0]  io_key,
  output [15:0] io_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] data [0:31]; // @[CAM.scala 22:17]
  wire [15:0] data_io_data_MPORT_data; // @[CAM.scala 22:17]
  wire [4:0] data_io_data_MPORT_addr; // @[CAM.scala 22:17]
  wire [15:0] data_MPORT_data; // @[CAM.scala 22:17]
  wire [4:0] data_MPORT_addr; // @[CAM.scala 22:17]
  wire  data_MPORT_mask; // @[CAM.scala 22:17]
  wire  data_MPORT_en; // @[CAM.scala 22:17]
  reg [31:0] free; // @[CAM.scala 21:21]
  wire [32:0] _free_sel_T = {free, 1'h0}; // @[package.scala 244:48]
  wire [31:0] _free_sel_T_2 = free | _free_sel_T[31:0]; // @[package.scala 244:43]
  wire [33:0] _free_sel_T_3 = {_free_sel_T_2, 2'h0}; // @[package.scala 244:48]
  wire [31:0] _free_sel_T_5 = _free_sel_T_2 | _free_sel_T_3[31:0]; // @[package.scala 244:43]
  wire [35:0] _free_sel_T_6 = {_free_sel_T_5, 4'h0}; // @[package.scala 244:48]
  wire [31:0] _free_sel_T_8 = _free_sel_T_5 | _free_sel_T_6[31:0]; // @[package.scala 244:43]
  wire [39:0] _free_sel_T_9 = {_free_sel_T_8, 8'h0}; // @[package.scala 244:48]
  wire [31:0] _free_sel_T_11 = _free_sel_T_8 | _free_sel_T_9[31:0]; // @[package.scala 244:43]
  wire [47:0] _free_sel_T_12 = {_free_sel_T_11, 16'h0}; // @[package.scala 244:48]
  wire [31:0] _free_sel_T_14 = _free_sel_T_11 | _free_sel_T_12[31:0]; // @[package.scala 244:43]
  wire [32:0] _free_sel_T_16 = {_free_sel_T_14, 1'h0}; // @[CAM.scala 24:39]
  wire [32:0] _free_sel_T_17 = ~_free_sel_T_16; // @[CAM.scala 24:18]
  wire [32:0] _GEN_5 = {{1'd0}, free}; // @[CAM.scala 24:45]
  wire [32:0] free_sel = _free_sel_T_17 & _GEN_5; // @[CAM.scala 24:45]
  wire [15:0] io_key_hi = free_sel[31:16]; // @[OneHot.scala 30:18]
  wire [15:0] io_key_lo = free_sel[15:0]; // @[OneHot.scala 31:18]
  wire  io_key_hi_1 = |io_key_hi; // @[OneHot.scala 32:14]
  wire [15:0] _io_key_T = io_key_hi | io_key_lo; // @[OneHot.scala 32:28]
  wire [7:0] io_key_hi_2 = _io_key_T[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] io_key_lo_1 = _io_key_T[7:0]; // @[OneHot.scala 31:18]
  wire  io_key_hi_3 = |io_key_hi_2; // @[OneHot.scala 32:14]
  wire [7:0] _io_key_T_1 = io_key_hi_2 | io_key_lo_1; // @[OneHot.scala 32:28]
  wire [3:0] io_key_hi_4 = _io_key_T_1[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] io_key_lo_2 = _io_key_T_1[3:0]; // @[OneHot.scala 31:18]
  wire  io_key_hi_5 = |io_key_hi_4; // @[OneHot.scala 32:14]
  wire [3:0] _io_key_T_2 = io_key_hi_4 | io_key_lo_2; // @[OneHot.scala 32:28]
  wire [1:0] io_key_hi_6 = _io_key_T_2[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] io_key_lo_3 = _io_key_T_2[1:0]; // @[OneHot.scala 31:18]
  wire  io_key_hi_7 = |io_key_hi_6; // @[OneHot.scala 32:14]
  wire [1:0] _io_key_T_3 = io_key_hi_6 | io_key_lo_3; // @[OneHot.scala 32:28]
  wire  io_key_lo_4 = _io_key_T_3[1]; // @[CircuitMath.scala 30:8]
  wire [3:0] io_key_lo_7 = {io_key_hi_3,io_key_hi_5,io_key_hi_7,io_key_lo_4}; // @[Cat.scala 30:58]
  wire  _T = io_alloc_ready & io_alloc_valid; // @[Decoupled.scala 40:37]
  wire  bypass = _T & 5'h0 == io_key; // @[CAM.scala 31:32]
  wire [32:0] clr = _T ? free_sel : 33'h0; // @[CAM.scala 35:16]
  wire [32:0] _free_T = ~clr; // @[CAM.scala 37:19]
  wire [32:0] _free_T_1 = _GEN_5 & _free_T; // @[CAM.scala 37:17]
  assign data_io_data_MPORT_addr = 5'h0;
  assign data_io_data_MPORT_data = data[data_io_data_MPORT_addr]; // @[CAM.scala 22:17]
  assign data_MPORT_data = io_alloc_bits;
  assign data_MPORT_addr = io_key;
  assign data_MPORT_mask = 1'h1;
  assign data_MPORT_en = io_alloc_ready & io_alloc_valid;
  assign io_alloc_ready = |free; // @[CAM.scala 27:26]
  assign io_key = {io_key_hi_1,io_key_lo_7}; // @[Cat.scala 30:58]
  assign io_data = bypass ? io_alloc_bits : data_io_data_MPORT_data; // @[CAM.scala 32:17]
  always @(posedge clock) begin
    if(data_MPORT_en & data_MPORT_mask) begin
      data[data_MPORT_addr] <= data_MPORT_data; // @[CAM.scala 22:17]
    end
    if (reset) begin // @[CAM.scala 21:21]
      free <= 32'hffffffff; // @[CAM.scala 21:21]
    end else begin
      free <= _free_T_1[31:0]; // @[CAM.scala 37:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    data[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  free = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SourceD(
  input         clock,
  input         reset,
  input         io_d_ready,
  output        io_d_valid,
  output [2:0]  io_d_bits_opcode,
  output [1:0]  io_d_bits_param,
  output [2:0]  io_d_bits_size,
  output [3:0]  io_d_bits_source,
  output [4:0]  io_d_bits_sink,
  output        io_d_bits_denied,
  output [31:0] io_d_bits_data,
  output        io_d_bits_corrupt,
  output        io_q_ready,
  input         io_q_valid,
  input  [31:0] io_q_bits,
  output [15:0] io_e_clSink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  cam_clock; // @[SourceD.scala 20:19]
  wire  cam_reset; // @[SourceD.scala 20:19]
  wire  cam_io_alloc_ready; // @[SourceD.scala 20:19]
  wire  cam_io_alloc_valid; // @[SourceD.scala 20:19]
  wire [15:0] cam_io_alloc_bits; // @[SourceD.scala 20:19]
  wire [4:0] cam_io_key; // @[SourceD.scala 20:19]
  wire [15:0] cam_io_data; // @[SourceD.scala 20:19]
  reg [1:0] state; // @[SourceD.scala 30:22]
  wire [2:0] opcode = io_q_bits[5:3]; // @[Parameters.scala 92:19]
  wire [2:0] param = io_q_bits[8:6]; // @[Parameters.scala 93:19]
  wire [3:0] size = io_q_bits[12:9]; // @[Parameters.scala 94:19]
  wire [2:0] domain = io_q_bits[15:13]; // @[Parameters.scala 95:19]
  wire [15:0] source = io_q_bits[31:16]; // @[Parameters.scala 96:19]
  wire  enable = state == 2'h0; // @[SourceD.scala 36:24]
  reg [2:0] r_1; // @[Reg.scala 15:16]
  wire [2:0] _GEN_1 = enable ? opcode : r_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [2:0] r_2; // @[Reg.scala 15:16]
  wire [2:0] _GEN_2 = enable ? param : r_2; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [3:0] r_3; // @[Reg.scala 15:16]
  wire [3:0] _GEN_3 = enable ? size : r_3; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [2:0] r_4; // @[Reg.scala 15:16]
  wire [2:0] _GEN_4 = enable ? domain : r_4; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [15:0] r_5; // @[Reg.scala 15:16]
  wire [15:0] _GEN_5 = enable ? source : r_5; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire  q_sink_enable = state == 2'h1; // @[SourceD.scala 36:24]
  reg [15:0] q_sink_r; // @[Reg.scala 15:16]
  wire  q_grant = _GEN_1 == 3'h4 | _GEN_1 == 3'h5; // @[SourceD.scala 47:47]
  reg [4:0] q_last_count; // @[Parameters.scala 126:24]
  wire [2:0] q_last_beats_beats_shiftAmount = size[2:0]; // @[OneHot.scala 64:49]
  wire [7:0] _q_last_beats_beats_T_1 = 8'h1 << q_last_beats_beats_shiftAmount; // @[OneHot.scala 65:12]
  wire [3:0] q_last_beats_beats_hi = _q_last_beats_beats_T_1[6:3]; // @[Parameters.scala 102:62]
  wire  q_last_beats_beats_lo = size <= 4'h2; // @[Parameters.scala 102:83]
  wire [4:0] q_last_beats_beats = {q_last_beats_beats_hi,q_last_beats_beats_lo}; // @[Cat.scala 30:58]
  wire  q_last_beats_grant = opcode == 3'h4 | opcode == 3'h5; // @[Parameters.scala 114:45]
  wire [4:0] _q_last_beats_c_T_1 = opcode[0] ? q_last_beats_beats : 5'h0; // @[Parameters.scala 118:16]
  wire [4:0] _GEN_40 = {{4'd0}, q_last_beats_grant}; // @[Parameters.scala 119:44]
  wire [4:0] q_last_beats_d = _q_last_beats_c_T_1 + _GEN_40; // @[Parameters.scala 119:44]
  wire  q_last_first = q_last_count == 5'h0; // @[Parameters.scala 128:23]
  wire  q_last = q_last_count == 5'h1 | q_last_first & q_last_beats_d == 5'h0; // @[Parameters.scala 129:35]
  wire  _q_last_T = io_q_ready & io_q_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _q_last_count_T_1 = q_last_count - 5'h1; // @[Parameters.scala 130:56]
  wire  _d_first_T = state != 2'h2; // @[SourceD.scala 49:33]
  reg  d_first; // @[Reg.scala 15:16]
  wire [1:0] s_maybe_data = q_last ? 2'h0 : 2'h2; // @[SourceD.scala 50:25]
  wire  _T_2 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_9 = _T_4 ? s_maybe_data : state; // @[Conditional.scala 39:67 SourceD.scala 56:31 SourceD.scala 30:22]
  wire  sink_ok = ~q_grant | cam_io_alloc_ready; // @[SourceD.scala 61:26]
  reg [4:0] sink_r; // @[Reg.scala 15:16]
  wire [4:0] _GEN_13 = d_first ? cam_io_key : sink_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire  stall = d_first & ~sink_ok; // @[SourceD.scala 63:23]
  wire  xmit = q_last | state == 2'h2; // @[SourceD.scala 64:22]
  wire [2:0] _GEN_15 = 3'h1 == _GEN_5[2:0] ? 3'h1 : 3'h0; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [2:0] _GEN_16 = 3'h2 == _GEN_5[2:0] ? 3'h2 : _GEN_15; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [2:0] _GEN_17 = 3'h3 == _GEN_5[2:0] ? 3'h3 : _GEN_16; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [2:0] _GEN_18 = 3'h4 == _GEN_5[2:0] ? 3'h4 : _GEN_17; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [2:0] _GEN_19 = 3'h5 == _GEN_5[2:0] ? 3'h5 : _GEN_18; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [2:0] _GEN_20 = 3'h6 == _GEN_5[2:0] ? 3'h6 : _GEN_19; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [2:0] _GEN_21 = 3'h7 == _GEN_5[2:0] ? 3'h7 : _GEN_20; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _GEN_23 = 3'h1 == _GEN_5[2:0] ? 4'h9 : 4'h8; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _GEN_24 = 3'h2 == _GEN_5[2:0] ? 4'ha : _GEN_23; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _GEN_25 = 3'h3 == _GEN_5[2:0] ? 4'hb : _GEN_24; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _GEN_26 = 3'h4 == _GEN_5[2:0] ? 4'hc : _GEN_25; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _GEN_27 = 3'h5 == _GEN_5[2:0] ? 4'hd : _GEN_26; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _GEN_28 = 3'h6 == _GEN_5[2:0] ? 4'he : _GEN_27; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _GEN_29 = 3'h7 == _GEN_5[2:0] ? 4'hf : _GEN_28; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _io_d_bits_source_WIRE_1 = {{1'd0}, _GEN_21}; // @[SourceD.scala 69:27 SourceD.scala 69:27]
  wire [3:0] _GEN_31 = 3'h1 == _GEN_4 ? _io_d_bits_source_WIRE_1 : 4'h0; // @[SourceD.scala 69:21 SourceD.scala 69:21]
  wire [3:0] _GEN_32 = 3'h2 == _GEN_4 ? _GEN_29 : _GEN_31; // @[SourceD.scala 69:21 SourceD.scala 69:21]
  wire [3:0] _GEN_33 = 3'h3 == _GEN_4 ? 4'h0 : _GEN_32; // @[SourceD.scala 69:21 SourceD.scala 69:21]
  wire [3:0] _GEN_34 = 3'h4 == _GEN_4 ? 4'h0 : _GEN_33; // @[SourceD.scala 69:21 SourceD.scala 69:21]
  wire [3:0] _GEN_35 = 3'h5 == _GEN_4 ? 4'h0 : _GEN_34; // @[SourceD.scala 69:21 SourceD.scala 69:21]
  wire [3:0] _GEN_36 = 3'h6 == _GEN_4 ? 4'h0 : _GEN_35; // @[SourceD.scala 69:21 SourceD.scala 69:21]
  wire  io_d_bits_corrupt_opdata = io_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  _io_d_valid_T = ~stall; // @[SourceD.scala 75:32]
  CAM_9 cam ( // @[SourceD.scala 20:19]
    .clock(cam_clock),
    .reset(cam_reset),
    .io_alloc_ready(cam_io_alloc_ready),
    .io_alloc_valid(cam_io_alloc_valid),
    .io_alloc_bits(cam_io_alloc_bits),
    .io_key(cam_io_key),
    .io_data(cam_io_data)
  );
  assign io_d_valid = io_q_valid & ~stall & xmit; // @[SourceD.scala 75:40]
  assign io_d_bits_opcode = enable ? opcode : r_1; // @[SourceD.scala 37:8]
  assign io_d_bits_param = _GEN_2[1:0]; // @[SourceD.scala 67:31]
  assign io_d_bits_size = _GEN_3[2:0]; // @[SourceD.scala 68:21]
  assign io_d_bits_source = 3'h7 == _GEN_4 ? 4'h0 : _GEN_36; // @[SourceD.scala 69:21 SourceD.scala 69:21]
  assign io_d_bits_sink = q_grant ? _GEN_13 : 5'h0; // @[SourceD.scala 70:27]
  assign io_d_bits_denied = _GEN_2[2]; // @[SourceD.scala 71:32]
  assign io_d_bits_data = io_q_bits; // @[SourceD.scala 72:21]
  assign io_d_bits_corrupt = io_d_bits_denied & io_d_bits_corrupt_opdata; // @[SourceD.scala 73:41]
  assign io_q_ready = io_d_ready & _io_d_valid_T | ~xmit; // @[SourceD.scala 76:40]
  assign io_e_clSink = cam_io_data; // @[SourceD.scala 82:15]
  assign cam_clock = clock;
  assign cam_reset = reset;
  assign cam_io_alloc_valid = q_grant & d_first & xmit & io_q_valid & io_d_ready; // @[SourceD.scala 78:66]
  assign cam_io_alloc_bits = q_sink_enable ? io_q_bits[15:0] : q_sink_r; // @[SourceD.scala 37:8]
  always @(posedge clock) begin
    if (reset) begin // @[SourceD.scala 30:22]
      state <= 2'h0; // @[SourceD.scala 30:22]
    end else if (_q_last_T) begin // @[SourceD.scala 52:22]
      if (_T_2) begin // @[Conditional.scala 40:58]
        if (q_grant) begin // @[SourceD.scala 54:37]
          state <= 2'h1;
        end else begin
          state <= s_maybe_data;
        end
      end else if (_T_3) begin // @[Conditional.scala 39:67]
        state <= s_maybe_data; // @[SourceD.scala 55:31]
      end else begin
        state <= _GEN_9;
      end
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_1 <= opcode; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_2 <= param; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_3 <= size; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_4 <= domain; // @[Reg.scala 16:23]
    end
    if (enable) begin // @[Reg.scala 16:19]
      r_5 <= source; // @[Reg.scala 16:23]
    end
    if (q_sink_enable) begin // @[Reg.scala 16:19]
      q_sink_r <= io_q_bits[15:0]; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Parameters.scala 126:24]
      q_last_count <= 5'h0; // @[Parameters.scala 126:24]
    end else if (_q_last_T) begin // @[Parameters.scala 130:21]
      if (q_last_first) begin // @[Parameters.scala 130:35]
        q_last_count <= q_last_beats_d;
      end else begin
        q_last_count <= _q_last_count_T_1;
      end
    end
    if (_q_last_T) begin // @[Reg.scala 16:19]
      d_first <= _d_first_T; // @[Reg.scala 16:23]
    end
    if (d_first) begin // @[Reg.scala 16:19]
      sink_r <= cam_io_key; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  r_4 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  r_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  q_sink_r = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  q_last_count = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  d_first = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sink_r = _RAND_9[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SourceE(
  input         io_e_ready,
  output        io_e_valid,
  output        io_e_bits_sink,
  output        io_q_ready,
  input         io_q_valid,
  input  [31:0] io_q_bits
);
  wire [15:0] q_sink = io_q_bits[31:16]; // @[Parameters.scala 96:19]
  assign io_e_valid = io_q_valid; // @[SourceE.scala 20:14]
  assign io_e_bits_sink = q_sink[0]; // @[SourceE.scala 21:18]
  assign io_q_ready = io_e_ready; // @[SourceE.scala 19:14]
endmodule
module HellaFlowQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] ram_R0_addr; // @[HellaQueue.scala 26:19]
  wire  ram_R0_en; // @[HellaQueue.scala 26:19]
  wire  ram_R0_clk; // @[HellaQueue.scala 26:19]
  wire [31:0] ram_R0_data; // @[HellaQueue.scala 26:19]
  wire [4:0] ram_W0_addr; // @[HellaQueue.scala 26:19]
  wire  ram_W0_en; // @[HellaQueue.scala 26:19]
  wire  ram_W0_clk; // @[HellaQueue.scala 26:19]
  wire [31:0] ram_W0_data; // @[HellaQueue.scala 26:19]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  reg [4:0] enq_ptr; // @[Counter.scala 60:40]
  reg [4:0] deq_ptr; // @[Counter.scala 60:40]
  wire  ptr_match = enq_ptr == deq_ptr; // @[HellaQueue.scala 20:27]
  reg  maybe_full; // @[HellaQueue.scala 15:23]
  wire  empty = ptr_match & ~maybe_full; // @[HellaQueue.scala 21:25]
  wire  do_flow = empty & io_deq_ready; // @[HellaQueue.scala 24:20]
  wire  _do_enq_T_1 = ~do_flow; // @[HellaQueue.scala 12:33]
  wire  do_enq = _do_enq_T & ~do_flow; // @[HellaQueue.scala 12:30]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = _do_deq_T & _do_enq_T_1; // @[HellaQueue.scala 13:30]
  wire [4:0] _enq_ptr_wrap_value_T_1 = enq_ptr + 5'h1; // @[Counter.scala 76:24]
  wire  wrap_wrap = deq_ptr == 5'h1f; // @[Counter.scala 72:24]
  wire [4:0] _wrap_value_T_1 = deq_ptr + 5'h1; // @[Counter.scala 76:24]
  wire  deq_done = do_deq & wrap_wrap; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire  full = ptr_match & maybe_full; // @[HellaQueue.scala 22:24]
  wire [4:0] _atLeastTwo_T_1 = enq_ptr - deq_ptr; // @[HellaQueue.scala 23:36]
  wire  atLeastTwo = full | _atLeastTwo_T_1 >= 5'h2; // @[HellaQueue.scala 23:25]
  wire [4:0] _raddr_T_2 = deq_done ? 5'h0 : _wrap_value_T_1; // @[HellaQueue.scala 32:36]
  reg  ram_out_valid; // @[HellaQueue.scala 33:26]
  ram ram ( // @[HellaQueue.scala 26:19]
    .R0_addr(ram_R0_addr),
    .R0_en(ram_R0_en),
    .R0_clk(ram_R0_clk),
    .R0_data(ram_R0_data),
    .W0_addr(ram_W0_addr),
    .W0_en(ram_W0_en),
    .W0_clk(ram_W0_clk),
    .W0_data(ram_W0_data)
  );
  assign io_enq_ready = ~full; // @[HellaQueue.scala 36:19]
  assign io_deq_valid = empty ? io_enq_valid : ram_out_valid; // @[HellaQueue.scala 35:22]
  assign io_deq_bits = empty ? io_enq_bits : ram_R0_data; // @[HellaQueue.scala 37:21]
  assign ram_R0_addr = io_deq_valid ? _raddr_T_2 : deq_ptr; // @[HellaQueue.scala 32:18]
  assign ram_R0_en = io_deq_ready & (atLeastTwo | ~io_deq_valid & ~empty); // @[HellaQueue.scala 31:26]
  assign ram_R0_clk = clock; // @[HellaQueue.scala 37:50 HellaQueue.scala 37:50]
  assign ram_W0_addr = enq_ptr; // @[HellaQueue.scala 27:17]
  assign ram_W0_en = _do_enq_T & ~do_flow; // @[HellaQueue.scala 12:30]
  assign ram_W0_clk = clock; // @[HellaQueue.scala 27:17]
  assign ram_W0_data = io_enq_bits; // @[HellaQueue.scala 27:17]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr <= 5'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Counter.scala 118:17]
      enq_ptr <= _enq_ptr_wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr <= 5'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Counter.scala 118:17]
      deq_ptr <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[HellaQueue.scala 15:23]
      maybe_full <= 1'h0; // @[HellaQueue.scala 15:23]
    end else if (do_enq != do_deq) begin // @[HellaQueue.scala 18:28]
      maybe_full <= do_enq; // @[HellaQueue.scala 18:41]
    end
    ram_out_valid <= io_deq_ready & (atLeastTwo | ~io_deq_valid & ~empty); // @[HellaQueue.scala 31:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_ptr = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  deq_ptr = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ram_out_valid = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:0]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign ram_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = 1'h0;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 254:25 Decoupled.scala 254:40 Decoupled.scala 241:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HellaQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
  wire  fq_clock; // @[HellaQueue.scala 43:18]
  wire  fq_reset; // @[HellaQueue.scala 43:18]
  wire  fq_io_enq_ready; // @[HellaQueue.scala 43:18]
  wire  fq_io_enq_valid; // @[HellaQueue.scala 43:18]
  wire [31:0] fq_io_enq_bits; // @[HellaQueue.scala 43:18]
  wire  fq_io_deq_ready; // @[HellaQueue.scala 43:18]
  wire  fq_io_deq_valid; // @[HellaQueue.scala 43:18]
  wire [31:0] fq_io_deq_bits; // @[HellaQueue.scala 43:18]
  wire  io_deq_q_clock; // @[Decoupled.scala 296:21]
  wire  io_deq_q_reset; // @[Decoupled.scala 296:21]
  wire  io_deq_q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  io_deq_q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] io_deq_q_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  io_deq_q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  io_deq_q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] io_deq_q_io_deq_bits; // @[Decoupled.scala 296:21]
  HellaFlowQueue fq ( // @[HellaQueue.scala 43:18]
    .clock(fq_clock),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits(fq_io_enq_bits),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits(fq_io_deq_bits)
  );
  Queue_6 io_deq_q ( // @[Decoupled.scala 296:21]
    .clock(io_deq_q_clock),
    .reset(io_deq_q_reset),
    .io_enq_ready(io_deq_q_io_enq_ready),
    .io_enq_valid(io_deq_q_io_enq_valid),
    .io_enq_bits(io_deq_q_io_enq_bits),
    .io_deq_ready(io_deq_q_io_deq_ready),
    .io_deq_valid(io_deq_q_io_deq_valid),
    .io_deq_bits(io_deq_q_io_deq_bits)
  );
  assign io_enq_ready = fq_io_enq_ready; // @[HellaQueue.scala 44:13]
  assign io_deq_valid = io_deq_q_io_deq_valid; // @[HellaQueue.scala 45:10]
  assign io_deq_bits = io_deq_q_io_deq_bits; // @[HellaQueue.scala 45:10]
  assign fq_clock = clock;
  assign fq_reset = reset;
  assign fq_io_enq_valid = io_enq_valid; // @[HellaQueue.scala 44:13]
  assign fq_io_enq_bits = io_enq_bits; // @[HellaQueue.scala 44:13]
  assign fq_io_deq_ready = io_deq_q_io_enq_ready; // @[Decoupled.scala 299:17]
  assign io_deq_q_clock = clock;
  assign io_deq_q_reset = reset;
  assign io_deq_q_io_enq_valid = fq_io_deq_valid; // @[Decoupled.scala 297:22]
  assign io_deq_q_io_enq_bits = fq_io_deq_bits; // @[Decoupled.scala 298:21]
  assign io_deq_q_io_deq_ready = io_deq_ready; // @[HellaQueue.scala 45:10]
endmodule
module AsyncResetSynchronizerPrimitiveShiftReg_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  sync_0; // @[SynchronizerReg.scala 51:87]
  reg  sync_1; // @[SynchronizerReg.scala 51:87]
  reg  sync_2; // @[SynchronizerReg.scala 51:87]
  assign io_q = sync_0; // @[SynchronizerReg.scala 59:8]
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      sync_0 <= 1'h0;
    end else begin
      sync_0 <= sync_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      sync_1 <= 1'h0;
    end else begin
      sync_1 <= sync_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      sync_2 <= 1'h0;
    end else begin
      sync_2 <= io_d;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sync_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sync_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    sync_0 = 1'h0;
  end
  if (reset) begin
    sync_1 = 1'h0;
  end
  if (reset) begin
    sync_2 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncResetSynchronizerShiftReg_w4_d3_i0(
  input        clock,
  input        reset,
  input  [3:0] io_d,
  output [3:0] io_q
);
  wire  output_chain_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_io_q; // @[ShiftReg.scala 45:23]
  wire  output_1 = output_chain_1_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire  output_0 = output_chain_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire [1:0] io_q_lo = {output_1,output_0}; // @[Cat.scala 30:58]
  wire  output_3 = output_chain_3_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire  output_2 = output_chain_2_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire [1:0] io_q_hi = {output_3,output_2}; // @[Cat.scala 30:58]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_clock),
    .reset(output_chain_reset),
    .io_d(output_chain_io_d),
    .io_q(output_chain_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_1 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_1_clock),
    .reset(output_chain_1_reset),
    .io_d(output_chain_1_io_d),
    .io_q(output_chain_1_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_2 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_2_clock),
    .reset(output_chain_2_reset),
    .io_d(output_chain_2_io_d),
    .io_q(output_chain_2_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_3 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_3_clock),
    .reset(output_chain_3_reset),
    .io_d(output_chain_3_io_d),
    .io_q(output_chain_3_io_q)
  );
  assign io_q = {io_q_hi,io_q_lo}; // @[Cat.scala 30:58]
  assign output_chain_clock = clock;
  assign output_chain_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_io_d = io_d[0]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_1_clock = clock;
  assign output_chain_1_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_1_io_d = io_d[1]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_2_clock = clock;
  assign output_chain_2_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_2_io_d = io_d[2]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_3_clock = clock;
  assign output_chain_3_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_3_io_d = io_d[3]; // @[SynchronizerReg.scala 87:41]
endmodule
module AsyncResetSynchronizerShiftReg_w1_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
  wire  output_chain_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_clock),
    .reset(output_chain_reset),
    .io_d(output_chain_io_d),
    .io_q(output_chain_io_q)
  );
  assign io_q = output_chain_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  assign output_chain_clock = clock;
  assign output_chain_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_io_d = io_d; // @[SynchronizerReg.scala 87:41]
endmodule
module AsyncValidSync(
  input   io_in,
  output  io_out,
  input   clock,
  input   reset
);
  wire  io_out_source_valid_0_clock; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_reset; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_io_d; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerShiftReg_w1_d3_i0 io_out_source_valid_0 ( // @[ShiftReg.scala 45:23]
    .clock(io_out_source_valid_0_clock),
    .reset(io_out_source_valid_0_reset),
    .io_d(io_out_source_valid_0_io_d),
    .io_q(io_out_source_valid_0_io_q)
  );
  assign io_out = io_out_source_valid_0_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  assign io_out_source_valid_0_clock = clock;
  assign io_out_source_valid_0_reset = reset;
  assign io_out_source_valid_0_io_d = io_in; // @[ShiftReg.scala 47:16]
endmodule
module AsyncQueueSource(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  output [31:0] io_async_mem_0,
  output [31:0] io_async_mem_1,
  output [31:0] io_async_mem_2,
  output [31:0] io_async_mem_3,
  output [31:0] io_async_mem_4,
  output [31:0] io_async_mem_5,
  output [31:0] io_async_mem_6,
  output [31:0] io_async_mem_7,
  input  [3:0]  io_async_ridx,
  output [3:0]  io_async_widx,
  input         io_async_safe_ridx_valid,
  output        io_async_safe_widx_valid,
  output        io_async_safe_source_reset_n,
  input         io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  ridx_ridx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  ridx_ridx_gray_reset; // @[ShiftReg.scala 45:23]
  wire [3:0] ridx_ridx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire [3:0] ridx_ridx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  source_valid_0_io_in; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_io_out; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_clock; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_reset; // @[AsyncQueue.scala 100:32]
  wire  source_valid_1_io_in; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_io_out; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_clock; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_reset; // @[AsyncQueue.scala 101:32]
  wire  sink_extend_io_in; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_io_out; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_clock; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_reset; // @[AsyncQueue.scala 103:30]
  wire  sink_valid_io_in; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_io_out; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_clock; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_reset; // @[AsyncQueue.scala 104:30]
  reg [31:0] mem_0; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_1; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_2; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_3; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_4; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_5; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_6; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_7; // @[AsyncQueue.scala 80:16]
  wire  _widx_T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  sink_ready = sink_valid_io_out;
  wire  _widx_T_2 = ~sink_ready; // @[AsyncQueue.scala 81:79]
  reg [3:0] widx_widx_bin; // @[AsyncQueue.scala 52:25]
  wire [3:0] _GEN_16 = {{3'd0}, _widx_T_1}; // @[AsyncQueue.scala 53:43]
  wire [3:0] _widx_incremented_T_1 = widx_widx_bin + _GEN_16; // @[AsyncQueue.scala 53:43]
  wire [3:0] widx_incremented = _widx_T_2 ? 4'h0 : _widx_incremented_T_1; // @[AsyncQueue.scala 53:23]
  wire [3:0] _GEN_17 = {{1'd0}, widx_incremented[3:1]}; // @[AsyncQueue.scala 54:17]
  wire [3:0] widx = widx_incremented ^ _GEN_17; // @[AsyncQueue.scala 54:17]
  wire [3:0] ridx = ridx_ridx_gray_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire [3:0] _ready_T = ridx ^ 4'hc; // @[AsyncQueue.scala 83:44]
  wire [2:0] _index_T_2 = {io_async_widx[3], 2'h0}; // @[AsyncQueue.scala 85:93]
  wire [2:0] index = io_async_widx[2:0] ^ _index_T_2; // @[AsyncQueue.scala 85:64]
  reg  ready_reg; // @[AsyncQueue.scala 88:56]
  reg [3:0] widx_gray; // @[AsyncQueue.scala 91:55]
  AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_ridx_gray ( // @[ShiftReg.scala 45:23]
    .clock(ridx_ridx_gray_clock),
    .reset(ridx_ridx_gray_reset),
    .io_d(ridx_ridx_gray_io_d),
    .io_q(ridx_ridx_gray_io_q)
  );
  AsyncValidSync source_valid_0 ( // @[AsyncQueue.scala 100:32]
    .io_in(source_valid_0_io_in),
    .io_out(source_valid_0_io_out),
    .clock(source_valid_0_clock),
    .reset(source_valid_0_reset)
  );
  AsyncValidSync source_valid_1 ( // @[AsyncQueue.scala 101:32]
    .io_in(source_valid_1_io_in),
    .io_out(source_valid_1_io_out),
    .clock(source_valid_1_clock),
    .reset(source_valid_1_reset)
  );
  AsyncValidSync sink_extend ( // @[AsyncQueue.scala 103:30]
    .io_in(sink_extend_io_in),
    .io_out(sink_extend_io_out),
    .clock(sink_extend_clock),
    .reset(sink_extend_reset)
  );
  AsyncValidSync sink_valid ( // @[AsyncQueue.scala 104:30]
    .io_in(sink_valid_io_in),
    .io_out(sink_valid_io_out),
    .clock(sink_valid_clock),
    .reset(sink_valid_reset)
  );
  assign io_enq_ready = ready_reg & sink_ready; // @[AsyncQueue.scala 89:29]
  assign io_async_mem_0 = mem_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1 = mem_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2 = mem_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3 = mem_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4 = mem_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5 = mem_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6 = mem_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7 = mem_7; // @[AsyncQueue.scala 96:31]
  assign io_async_widx = widx_gray; // @[AsyncQueue.scala 92:17]
  assign io_async_safe_widx_valid = source_valid_1_io_out; // @[AsyncQueue.scala 117:20]
  assign io_async_safe_source_reset_n = ~reset; // @[AsyncQueue.scala 121:27]
  assign ridx_ridx_gray_clock = clock;
  assign ridx_ridx_gray_reset = reset;
  assign ridx_ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 47:16]
  assign source_valid_0_io_in = 1'h1; // @[AsyncQueue.scala 115:26]
  assign source_valid_0_clock = clock; // @[AsyncQueue.scala 110:26]
  assign source_valid_0_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 105:65]
  assign source_valid_1_io_in = source_valid_0_io_out; // @[AsyncQueue.scala 116:26]
  assign source_valid_1_clock = clock; // @[AsyncQueue.scala 111:26]
  assign source_valid_1_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 106:65]
  assign sink_extend_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 118:23]
  assign sink_extend_clock = clock; // @[AsyncQueue.scala 112:26]
  assign sink_extend_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 107:65]
  assign sink_valid_io_in = sink_extend_io_out; // @[AsyncQueue.scala 119:22]
  assign sink_valid_clock = clock; // @[AsyncQueue.scala 113:26]
  assign sink_valid_reset = reset; // @[AsyncQueue.scala 108:35]
  always @(posedge clock) begin
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h0 == index) begin // @[AsyncQueue.scala 86:37]
        mem_0 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h1 == index) begin // @[AsyncQueue.scala 86:37]
        mem_1 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h2 == index) begin // @[AsyncQueue.scala 86:37]
        mem_2 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h3 == index) begin // @[AsyncQueue.scala 86:37]
        mem_3 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h4 == index) begin // @[AsyncQueue.scala 86:37]
        mem_4 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h5 == index) begin // @[AsyncQueue.scala 86:37]
        mem_5 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h6 == index) begin // @[AsyncQueue.scala 86:37]
        mem_6 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h7 == index) begin // @[AsyncQueue.scala 86:37]
        mem_7 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      widx_widx_bin <= 4'h0;
    end else if (_widx_T_2) begin
      widx_widx_bin <= 4'h0;
    end else begin
      widx_widx_bin <= _widx_incremented_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ready_reg <= 1'h0;
    end else begin
      ready_reg <= sink_ready & widx != _ready_T;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      widx_gray <= 4'h0;
    end else begin
      widx_gray <= widx_incremented ^ _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  widx_widx_bin = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  ready_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  widx_gray = _RAND_10[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    widx_widx_bin = 4'h0;
  end
  if (reset) begin
    ready_reg = 1'h0;
  end
  if (reset) begin
    widx_gray = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncResetSynchronizerShiftReg_w1_d3_i0_20(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
  wire  output_chain_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_clock),
    .reset(output_chain_reset),
    .io_d(output_chain_io_d),
    .io_q(output_chain_io_q)
  );
  assign io_q = output_chain_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  assign output_chain_clock = clock;
  assign output_chain_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_io_d = io_d; // @[SynchronizerReg.scala 87:41]
endmodule
module AsyncQueueSource_5(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input  [19:0] io_enq_bits_a,
  input  [19:0] io_enq_bits_b,
  input  [19:0] io_enq_bits_c,
  input  [19:0] io_enq_bits_d,
  input  [19:0] io_enq_bits_e,
  output [19:0] io_async_mem_0_a,
  output [19:0] io_async_mem_0_b,
  output [19:0] io_async_mem_0_c,
  output [19:0] io_async_mem_0_d,
  output [19:0] io_async_mem_0_e,
  input         io_async_ridx,
  output        io_async_widx,
  input         io_async_safe_ridx_valid,
  output        io_async_safe_widx_valid,
  output        io_async_safe_source_reset_n,
  input         io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  ridx_ridx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  ridx_ridx_gray_reset; // @[ShiftReg.scala 45:23]
  wire  ridx_ridx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire  ridx_ridx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  source_valid_0_io_in; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_io_out; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_clock; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_reset; // @[AsyncQueue.scala 100:32]
  wire  source_valid_1_io_in; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_io_out; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_clock; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_reset; // @[AsyncQueue.scala 101:32]
  wire  sink_extend_io_in; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_io_out; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_clock; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_reset; // @[AsyncQueue.scala 103:30]
  wire  sink_valid_io_in; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_io_out; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_clock; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_reset; // @[AsyncQueue.scala 104:30]
  reg [19:0] mem_0_a; // @[AsyncQueue.scala 80:16]
  reg [19:0] mem_0_b; // @[AsyncQueue.scala 80:16]
  reg [19:0] mem_0_c; // @[AsyncQueue.scala 80:16]
  reg [19:0] mem_0_d; // @[AsyncQueue.scala 80:16]
  reg [19:0] mem_0_e; // @[AsyncQueue.scala 80:16]
  wire  sink_ready = sink_valid_io_out;
  wire  _widx_T_2 = ~sink_ready; // @[AsyncQueue.scala 81:79]
  reg  widx_widx_bin; // @[AsyncQueue.scala 52:25]
  wire  widx_incremented = _widx_T_2 ? 1'h0 : widx_widx_bin + io_enq_ready; // @[AsyncQueue.scala 53:23]
  wire  ridx = ridx_ridx_gray_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  reg  ready_reg; // @[AsyncQueue.scala 88:56]
  reg  widx_gray; // @[AsyncQueue.scala 91:55]
  AsyncResetSynchronizerShiftReg_w1_d3_i0_20 ridx_ridx_gray ( // @[ShiftReg.scala 45:23]
    .clock(ridx_ridx_gray_clock),
    .reset(ridx_ridx_gray_reset),
    .io_d(ridx_ridx_gray_io_d),
    .io_q(ridx_ridx_gray_io_q)
  );
  AsyncValidSync source_valid_0 ( // @[AsyncQueue.scala 100:32]
    .io_in(source_valid_0_io_in),
    .io_out(source_valid_0_io_out),
    .clock(source_valid_0_clock),
    .reset(source_valid_0_reset)
  );
  AsyncValidSync source_valid_1 ( // @[AsyncQueue.scala 101:32]
    .io_in(source_valid_1_io_in),
    .io_out(source_valid_1_io_out),
    .clock(source_valid_1_clock),
    .reset(source_valid_1_reset)
  );
  AsyncValidSync sink_extend ( // @[AsyncQueue.scala 103:30]
    .io_in(sink_extend_io_in),
    .io_out(sink_extend_io_out),
    .clock(sink_extend_clock),
    .reset(sink_extend_reset)
  );
  AsyncValidSync sink_valid ( // @[AsyncQueue.scala 104:30]
    .io_in(sink_valid_io_in),
    .io_out(sink_valid_io_out),
    .clock(sink_valid_clock),
    .reset(sink_valid_reset)
  );
  assign io_enq_ready = ready_reg & sink_ready; // @[AsyncQueue.scala 89:29]
  assign io_async_mem_0_a = mem_0_a; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_b = mem_0_b; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_c = mem_0_c; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_d = mem_0_d; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_e = mem_0_e; // @[AsyncQueue.scala 96:31]
  assign io_async_widx = widx_gray; // @[AsyncQueue.scala 92:17]
  assign io_async_safe_widx_valid = source_valid_1_io_out; // @[AsyncQueue.scala 117:20]
  assign io_async_safe_source_reset_n = ~reset; // @[AsyncQueue.scala 121:27]
  assign ridx_ridx_gray_clock = clock;
  assign ridx_ridx_gray_reset = reset;
  assign ridx_ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 47:16]
  assign source_valid_0_io_in = 1'h1; // @[AsyncQueue.scala 115:26]
  assign source_valid_0_clock = clock; // @[AsyncQueue.scala 110:26]
  assign source_valid_0_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 105:65]
  assign source_valid_1_io_in = source_valid_0_io_out; // @[AsyncQueue.scala 116:26]
  assign source_valid_1_clock = clock; // @[AsyncQueue.scala 111:26]
  assign source_valid_1_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 106:65]
  assign sink_extend_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 118:23]
  assign sink_extend_clock = clock; // @[AsyncQueue.scala 112:26]
  assign sink_extend_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 107:65]
  assign sink_valid_io_in = sink_extend_io_out; // @[AsyncQueue.scala 119:22]
  assign sink_valid_clock = clock; // @[AsyncQueue.scala 113:26]
  assign sink_valid_reset = reset; // @[AsyncQueue.scala 108:35]
  always @(posedge clock) begin
    if (io_enq_ready) begin // @[AsyncQueue.scala 86:24]
      mem_0_a <= io_enq_bits_a; // @[AsyncQueue.scala 86:37]
    end
    if (io_enq_ready) begin // @[AsyncQueue.scala 86:24]
      mem_0_b <= io_enq_bits_b; // @[AsyncQueue.scala 86:37]
    end
    if (io_enq_ready) begin // @[AsyncQueue.scala 86:24]
      mem_0_c <= io_enq_bits_c; // @[AsyncQueue.scala 86:37]
    end
    if (io_enq_ready) begin // @[AsyncQueue.scala 86:24]
      mem_0_d <= io_enq_bits_d; // @[AsyncQueue.scala 86:37]
    end
    if (io_enq_ready) begin // @[AsyncQueue.scala 86:24]
      mem_0_e <= io_enq_bits_e; // @[AsyncQueue.scala 86:37]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      widx_widx_bin <= 1'h0;
    end else if (_widx_T_2) begin
      widx_widx_bin <= 1'h0;
    end else begin
      widx_widx_bin <= widx_widx_bin + io_enq_ready;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ready_reg <= 1'h0;
    end else begin
      ready_reg <= sink_ready & widx_incremented != (ridx ^ 1'h1);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      widx_gray <= 1'h0;
    end else if (_widx_T_2) begin
      widx_gray <= 1'h0;
    end else begin
      widx_gray <= widx_widx_bin + io_enq_ready;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_a = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_b = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  mem_0_c = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  mem_0_d = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  mem_0_e = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  widx_widx_bin = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ready_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  widx_gray = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    widx_widx_bin = 1'h0;
  end
  if (reset) begin
    ready_reg = 1'h0;
  end
  if (reset) begin
    widx_gray = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RX(
  input         clock,
  input         reset,
  input         io_b2c_send,
  input  [7:0]  io_b2c_data,
  output [31:0] io_a_mem_0,
  output [31:0] io_a_mem_1,
  output [31:0] io_a_mem_2,
  output [31:0] io_a_mem_3,
  output [31:0] io_a_mem_4,
  output [31:0] io_a_mem_5,
  output [31:0] io_a_mem_6,
  output [31:0] io_a_mem_7,
  input  [3:0]  io_a_ridx,
  output [3:0]  io_a_widx,
  input         io_a_safe_ridx_valid,
  output        io_a_safe_widx_valid,
  output        io_a_safe_source_reset_n,
  input         io_a_safe_sink_reset_n,
  output [31:0] io_bmem_0,
  output [31:0] io_bmem_1,
  output [31:0] io_bmem_2,
  output [31:0] io_bmem_3,
  output [31:0] io_bmem_4,
  output [31:0] io_bmem_5,
  output [31:0] io_bmem_6,
  output [31:0] io_bmem_7,
  input  [3:0]  io_bridx,
  output [3:0]  io_bwidx,
  input         io_bsafe_ridx_valid,
  output        io_bsafe_widx_valid,
  output        io_bsafe_source_reset_n,
  input         io_bsafe_sink_reset_n,
  output [31:0] io_c_mem_0,
  output [31:0] io_c_mem_1,
  output [31:0] io_c_mem_2,
  output [31:0] io_c_mem_3,
  output [31:0] io_c_mem_4,
  output [31:0] io_c_mem_5,
  output [31:0] io_c_mem_6,
  output [31:0] io_c_mem_7,
  input  [3:0]  io_c_ridx,
  output [3:0]  io_c_widx,
  input         io_c_safe_ridx_valid,
  output        io_c_safe_widx_valid,
  output        io_c_safe_source_reset_n,
  input         io_c_safe_sink_reset_n,
  output [31:0] io_d_mem_0,
  output [31:0] io_d_mem_1,
  output [31:0] io_d_mem_2,
  output [31:0] io_d_mem_3,
  output [31:0] io_d_mem_4,
  output [31:0] io_d_mem_5,
  output [31:0] io_d_mem_6,
  output [31:0] io_d_mem_7,
  input  [3:0]  io_d_ridx,
  output [3:0]  io_d_widx,
  input         io_d_safe_ridx_valid,
  output        io_d_safe_widx_valid,
  output        io_d_safe_source_reset_n,
  input         io_d_safe_sink_reset_n,
  output [31:0] io_e_mem_0,
  output [31:0] io_e_mem_1,
  output [31:0] io_e_mem_2,
  output [31:0] io_e_mem_3,
  output [31:0] io_e_mem_4,
  output [31:0] io_e_mem_5,
  output [31:0] io_e_mem_6,
  output [31:0] io_e_mem_7,
  input  [3:0]  io_e_ridx,
  output [3:0]  io_e_widx,
  input         io_e_safe_ridx_valid,
  output        io_e_safe_widx_valid,
  output        io_e_safe_source_reset_n,
  input         io_e_safe_sink_reset_n,
  output [19:0] io_rxc_mem_0_a,
  output [19:0] io_rxc_mem_0_b,
  output [19:0] io_rxc_mem_0_c,
  output [19:0] io_rxc_mem_0_d,
  output [19:0] io_rxc_mem_0_e,
  input         io_rxc_ridx,
  output        io_rxc_widx,
  input         io_rxc_safe_ridx_valid,
  output        io_rxc_safe_widx_valid,
  output        io_rxc_safe_source_reset_n,
  input         io_rxc_safe_sink_reset_n,
  output [19:0] io_txc_mem_0_a,
  output [19:0] io_txc_mem_0_b,
  output [19:0] io_txc_mem_0_c,
  output [19:0] io_txc_mem_0_d,
  output [19:0] io_txc_mem_0_e,
  input         io_txc_ridx,
  output        io_txc_widx,
  input         io_txc_safe_ridx_valid,
  output        io_txc_safe_widx_valid,
  output        io_txc_safe_source_reset_n,
  input         io_txc_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  hqa_clock; // @[RX.scala 50:19]
  wire  hqa_reset; // @[RX.scala 50:19]
  wire  hqa_io_enq_ready; // @[RX.scala 50:19]
  wire  hqa_io_enq_valid; // @[RX.scala 50:19]
  wire [31:0] hqa_io_enq_bits; // @[RX.scala 50:19]
  wire  hqa_io_deq_ready; // @[RX.scala 50:19]
  wire  hqa_io_deq_valid; // @[RX.scala 50:19]
  wire [31:0] hqa_io_deq_bits; // @[RX.scala 50:19]
  wire  hqb_clock; // @[RX.scala 51:19]
  wire  hqb_reset; // @[RX.scala 51:19]
  wire  hqb_io_enq_ready; // @[RX.scala 51:19]
  wire  hqb_io_enq_valid; // @[RX.scala 51:19]
  wire [31:0] hqb_io_enq_bits; // @[RX.scala 51:19]
  wire  hqb_io_deq_ready; // @[RX.scala 51:19]
  wire  hqb_io_deq_valid; // @[RX.scala 51:19]
  wire [31:0] hqb_io_deq_bits; // @[RX.scala 51:19]
  wire  hqc_clock; // @[RX.scala 52:19]
  wire  hqc_reset; // @[RX.scala 52:19]
  wire  hqc_io_enq_ready; // @[RX.scala 52:19]
  wire  hqc_io_enq_valid; // @[RX.scala 52:19]
  wire [31:0] hqc_io_enq_bits; // @[RX.scala 52:19]
  wire  hqc_io_deq_ready; // @[RX.scala 52:19]
  wire  hqc_io_deq_valid; // @[RX.scala 52:19]
  wire [31:0] hqc_io_deq_bits; // @[RX.scala 52:19]
  wire  hqd_clock; // @[RX.scala 53:19]
  wire  hqd_reset; // @[RX.scala 53:19]
  wire  hqd_io_enq_ready; // @[RX.scala 53:19]
  wire  hqd_io_enq_valid; // @[RX.scala 53:19]
  wire [31:0] hqd_io_enq_bits; // @[RX.scala 53:19]
  wire  hqd_io_deq_ready; // @[RX.scala 53:19]
  wire  hqd_io_deq_valid; // @[RX.scala 53:19]
  wire [31:0] hqd_io_deq_bits; // @[RX.scala 53:19]
  wire  hqe_clock; // @[RX.scala 54:19]
  wire  hqe_reset; // @[RX.scala 54:19]
  wire  hqe_io_enq_ready; // @[RX.scala 54:19]
  wire  hqe_io_enq_valid; // @[RX.scala 54:19]
  wire [31:0] hqe_io_enq_bits; // @[RX.scala 54:19]
  wire  hqe_io_deq_ready; // @[RX.scala 54:19]
  wire  hqe_io_deq_valid; // @[RX.scala 54:19]
  wire [31:0] hqe_io_deq_bits; // @[RX.scala 54:19]
  wire  io_a_source_clock; // @[AsyncQueue.scala 216:24]
  wire  io_a_source_reset; // @[AsyncQueue.scala 216:24]
  wire  io_a_source_io_enq_ready; // @[AsyncQueue.scala 216:24]
  wire  io_a_source_io_enq_valid; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_enq_bits; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_async_mem_0; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_async_mem_1; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_async_mem_2; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_async_mem_3; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_async_mem_4; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_async_mem_5; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_async_mem_6; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_a_source_io_async_mem_7; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_a_source_io_async_ridx; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_a_source_io_async_widx; // @[AsyncQueue.scala 216:24]
  wire  io_a_source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_a_source_io_async_safe_widx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_a_source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_a_source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_bsource_clock; // @[AsyncQueue.scala 216:24]
  wire  io_bsource_reset; // @[AsyncQueue.scala 216:24]
  wire  io_bsource_io_enq_ready; // @[AsyncQueue.scala 216:24]
  wire  io_bsource_io_enq_valid; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_enq_bits; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_async_mem_0; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_async_mem_1; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_async_mem_2; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_async_mem_3; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_async_mem_4; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_async_mem_5; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_async_mem_6; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_bsource_io_async_mem_7; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_bsource_io_async_ridx; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_bsource_io_async_widx; // @[AsyncQueue.scala 216:24]
  wire  io_bsource_io_async_safe_ridx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_bsource_io_async_safe_widx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_bsource_io_async_safe_source_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_bsource_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_c_source_clock; // @[AsyncQueue.scala 216:24]
  wire  io_c_source_reset; // @[AsyncQueue.scala 216:24]
  wire  io_c_source_io_enq_ready; // @[AsyncQueue.scala 216:24]
  wire  io_c_source_io_enq_valid; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_enq_bits; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_async_mem_0; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_async_mem_1; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_async_mem_2; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_async_mem_3; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_async_mem_4; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_async_mem_5; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_async_mem_6; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_c_source_io_async_mem_7; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_c_source_io_async_ridx; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_c_source_io_async_widx; // @[AsyncQueue.scala 216:24]
  wire  io_c_source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_c_source_io_async_safe_widx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_c_source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_c_source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_d_source_clock; // @[AsyncQueue.scala 216:24]
  wire  io_d_source_reset; // @[AsyncQueue.scala 216:24]
  wire  io_d_source_io_enq_ready; // @[AsyncQueue.scala 216:24]
  wire  io_d_source_io_enq_valid; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_enq_bits; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_async_mem_0; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_async_mem_1; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_async_mem_2; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_async_mem_3; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_async_mem_4; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_async_mem_5; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_async_mem_6; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_d_source_io_async_mem_7; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_d_source_io_async_ridx; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_d_source_io_async_widx; // @[AsyncQueue.scala 216:24]
  wire  io_d_source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_d_source_io_async_safe_widx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_d_source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_d_source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_e_source_clock; // @[AsyncQueue.scala 216:24]
  wire  io_e_source_reset; // @[AsyncQueue.scala 216:24]
  wire  io_e_source_io_enq_ready; // @[AsyncQueue.scala 216:24]
  wire  io_e_source_io_enq_valid; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_enq_bits; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_async_mem_0; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_async_mem_1; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_async_mem_2; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_async_mem_3; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_async_mem_4; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_async_mem_5; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_async_mem_6; // @[AsyncQueue.scala 216:24]
  wire [31:0] io_e_source_io_async_mem_7; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_e_source_io_async_ridx; // @[AsyncQueue.scala 216:24]
  wire [3:0] io_e_source_io_async_widx; // @[AsyncQueue.scala 216:24]
  wire  io_e_source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_e_source_io_async_safe_widx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_e_source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_e_source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_clock; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_reset; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_io_enq_ready; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_enq_bits_a; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_enq_bits_b; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_enq_bits_c; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_enq_bits_d; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_enq_bits_e; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_async_mem_0_a; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_async_mem_0_b; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_async_mem_0_c; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_async_mem_0_d; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_txc_source_io_async_mem_0_e; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_io_async_ridx; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_io_async_widx; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_io_async_safe_widx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_txc_source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_clock; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_reset; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_io_enq_ready; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_enq_bits_a; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_enq_bits_b; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_enq_bits_c; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_enq_bits_d; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_enq_bits_e; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_async_mem_0_a; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_async_mem_0_b; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_async_mem_0_c; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_async_mem_0_d; // @[AsyncQueue.scala 216:24]
  wire [19:0] io_rxc_source_io_async_mem_0_e; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_io_async_ridx; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_io_async_widx; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_io_async_safe_widx_valid; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 216:24]
  wire  io_rxc_source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 216:24]
  reg [7:0] b2c_data_REG; // @[RX.scala 24:33]
  reg [7:0] b2c_data; // @[RX.scala 24:25]
  reg  b2c_send_REG; // @[RX.scala 25:33]
  reg  b2c_send; // @[RX.scala 25:25]
  reg [1:0] beatCnt; // @[RX.scala 27:24]
  reg [31:0] b2c_data_concat; // @[RX.scala 28:32]
  reg  b2c_data_valid; // @[RX.scala 29:31]
  wire [1:0] _beatCnt_T_1 = beatCnt + 2'h1; // @[RX.scala 31:24]
  wire [39:0] _GEN_20 = {b2c_data_concat, 8'h0}; // @[RX.scala 32:41]
  wire [46:0] _b2c_data_concat_T = {{7'd0}, _GEN_20}; // @[RX.scala 32:41]
  wire [46:0] _GEN_21 = {{39'd0}, b2c_data}; // @[RX.scala 32:49]
  wire [46:0] _b2c_data_concat_T_1 = _b2c_data_concat_T | _GEN_21; // @[RX.scala 32:49]
  wire [46:0] _GEN_1 = b2c_send ? _b2c_data_concat_T_1 : {{15'd0}, b2c_data_concat}; // @[RX.scala 30:18 RX.scala 32:21 RX.scala 28:32]
  reg [4:0] first_count; // @[Parameters.scala 126:24]
  wire [2:0] first_beats_format = b2c_data_concat[2:0]; // @[Parameters.scala 91:19]
  wire [2:0] first_beats_opcode = b2c_data_concat[5:3]; // @[Parameters.scala 92:19]
  wire [3:0] first_beats_size = b2c_data_concat[12:9]; // @[Parameters.scala 94:19]
  wire [2:0] first_beats_beats_shiftAmount = first_beats_size[2:0]; // @[OneHot.scala 64:49]
  wire [7:0] _first_beats_beats_T_1 = 8'h1 << first_beats_beats_shiftAmount; // @[OneHot.scala 65:12]
  wire [3:0] first_beats_beats_hi = _first_beats_beats_T_1[6:3]; // @[Parameters.scala 102:62]
  wire  first_beats_beats_lo = first_beats_size <= 4'h2; // @[Parameters.scala 102:83]
  wire [4:0] first_beats_beats = {first_beats_beats_hi,first_beats_beats_lo}; // @[Cat.scala 30:58]
  wire  first_beats_masks_hi = _first_beats_beats_T_1[6]; // @[Parameters.scala 107:62]
  wire  first_beats_masks_lo = first_beats_size <= 4'h5; // @[Parameters.scala 107:83]
  wire [1:0] first_beats_masks = {first_beats_masks_hi,first_beats_masks_lo}; // @[Cat.scala 30:58]
  wire  first_beats_grant = first_beats_opcode == 3'h4 | first_beats_opcode == 3'h5; // @[Parameters.scala 114:45]
  wire  first_beats_partial = first_beats_opcode == 3'h1; // @[Parameters.scala 115:26]
  wire [4:0] _first_beats_a_T_1 = first_beats_opcode[2] ? 5'h0 : first_beats_beats; // @[Parameters.scala 116:16]
  wire [4:0] _first_beats_a_T_3 = _first_beats_a_T_1 + 5'h2; // @[Parameters.scala 116:44]
  wire [1:0] _first_beats_a_T_4 = first_beats_partial ? first_beats_masks : 2'h0; // @[Parameters.scala 116:59]
  wire [4:0] _GEN_22 = {{3'd0}, _first_beats_a_T_4}; // @[Parameters.scala 116:54]
  wire [4:0] first_beats_a = _first_beats_a_T_3 + _GEN_22; // @[Parameters.scala 116:54]
  wire [4:0] _first_beats_c_T_1 = first_beats_opcode[0] ? first_beats_beats : 5'h0; // @[Parameters.scala 118:16]
  wire [4:0] first_beats_c = _first_beats_c_T_1 + 5'h2; // @[Parameters.scala 118:44]
  wire [4:0] _GEN_24 = {{4'd0}, first_beats_grant}; // @[Parameters.scala 119:44]
  wire [4:0] first_beats_d = _first_beats_c_T_1 + _GEN_24; // @[Parameters.scala 119:44]
  wire  first = first_count == 5'h0; // @[Parameters.scala 128:23]
  wire [4:0] _GEN_3 = 3'h1 == first_beats_format ? first_beats_a : first_beats_a; // @[Parameters.scala 129:54 Parameters.scala 129:54]
  wire [4:0] _GEN_4 = 3'h2 == first_beats_format ? first_beats_c : _GEN_3; // @[Parameters.scala 129:54 Parameters.scala 129:54]
  wire [4:0] _GEN_5 = 3'h3 == first_beats_format ? first_beats_d : _GEN_4; // @[Parameters.scala 129:54 Parameters.scala 129:54]
  wire [4:0] _GEN_6 = 3'h4 == first_beats_format ? 5'h0 : _GEN_5; // @[Parameters.scala 129:54 Parameters.scala 129:54]
  wire [4:0] _first_count_T_1 = first_count - 5'h1; // @[Parameters.scala 130:56]
  wire  formatValid = b2c_data_valid & first; // @[RX.scala 45:33]
  reg [2:0] format_r; // @[Reg.scala 15:16]
  wire [2:0] _GEN_9 = formatValid ? first_beats_format : format_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire [7:0] formatOH = 8'h1 << _GEN_9; // @[OneHot.scala 58:35]
  reg [19:0] tx_a; // @[RX.scala 73:19]
  reg [19:0] tx_b; // @[RX.scala 73:19]
  reg [19:0] tx_c; // @[RX.scala 73:19]
  reg [19:0] tx_d; // @[RX.scala 73:19]
  reg [19:0] tx_e; // @[RX.scala 73:19]
  reg [19:0] rx_a; // @[RX.scala 74:19]
  reg [19:0] rx_b; // @[RX.scala 74:19]
  reg [19:0] rx_c; // @[RX.scala 74:19]
  reg [19:0] rx_d; // @[RX.scala 74:19]
  reg [19:0] rx_e; // @[RX.scala 74:19]
  wire  _rxInc_a_T = hqa_io_deq_ready & hqa_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _rxInc_bT = hqb_io_deq_ready & hqb_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _rxInc_c_T = hqc_io_deq_ready & hqc_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _rxInc_d_T = hqd_io_deq_ready & hqd_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _rxInc_e_T = hqe_io_deq_ready & hqe_io_deq_valid; // @[Decoupled.scala 40:37]
  wire [4:0] txInc_out_a_shiftAmount = b2c_data_concat[11:7]; // @[Bundles.scala 87:28]
  wire [31:0] _txInc_out_a_T_3 = 32'h1 << txInc_out_a_shiftAmount; // @[OneHot.scala 65:12]
  wire [19:0] txInc_out_a = txInc_out_a_shiftAmount > 5'h14 ? 20'hfffff : _txInc_out_a_T_3[20:1]; // @[Bundles.scala 83:10]
  wire [4:0] txInc_out_bshiftAmount = b2c_data_concat[16:12]; // @[Bundles.scala 88:28]
  wire [31:0] _txInc_out_bT_3 = 32'h1 << txInc_out_bshiftAmount; // @[OneHot.scala 65:12]
  wire [19:0] txInc_out_b = txInc_out_bshiftAmount > 5'h14 ? 20'hfffff : _txInc_out_bT_3[20:1]; // @[Bundles.scala 83:10]
  wire [4:0] txInc_out_c_shiftAmount = b2c_data_concat[21:17]; // @[Bundles.scala 89:28]
  wire [31:0] _txInc_out_c_T_3 = 32'h1 << txInc_out_c_shiftAmount; // @[OneHot.scala 65:12]
  wire [19:0] txInc_out_c = txInc_out_c_shiftAmount > 5'h14 ? 20'hfffff : _txInc_out_c_T_3[20:1]; // @[Bundles.scala 83:10]
  wire [4:0] txInc_out_d_shiftAmount = b2c_data_concat[26:22]; // @[Bundles.scala 90:28]
  wire [31:0] _txInc_out_d_T_3 = 32'h1 << txInc_out_d_shiftAmount; // @[OneHot.scala 65:12]
  wire [19:0] txInc_out_d = txInc_out_d_shiftAmount > 5'h14 ? 20'hfffff : _txInc_out_d_T_3[20:1]; // @[Bundles.scala 83:10]
  wire [4:0] txInc_out_e_shiftAmount = b2c_data_concat[31:27]; // @[Bundles.scala 91:28]
  wire [31:0] _txInc_out_e_T_3 = 32'h1 << txInc_out_e_shiftAmount; // @[OneHot.scala 65:12]
  wire [19:0] txInc_out_e = txInc_out_e_shiftAmount > 5'h14 ? 20'hfffff : _txInc_out_e_T_3[20:1]; // @[Bundles.scala 83:10]
  wire [19:0] txInc_a = b2c_data_valid & formatOH[5] ? txInc_out_a : 20'h0; // @[RX.scala 93:18]
  wire [19:0] txInc_b = b2c_data_valid & formatOH[5] ? txInc_out_b : 20'h0; // @[RX.scala 93:18]
  wire [19:0] txInc_c = b2c_data_valid & formatOH[5] ? txInc_out_c : 20'h0; // @[RX.scala 93:18]
  wire [19:0] txInc_d = b2c_data_valid & formatOH[5] ? txInc_out_d : 20'h0; // @[RX.scala 93:18]
  wire [19:0] txInc_e = b2c_data_valid & formatOH[5] ? txInc_out_e : 20'h0; // @[RX.scala 93:18]
  wire [20:0] tx_z = tx_a + txInc_a; // @[Bundles.scala 38:17]
  wire [20:0] _tx_out_a_T_3 = |tx_z[20] ? 21'hfffff : tx_z; // @[Bundles.scala 39:15]
  wire [20:0] tx_z_1 = tx_b + txInc_b; // @[Bundles.scala 38:17]
  wire [20:0] _tx_out_bT_3 = |tx_z_1[20] ? 21'hfffff : tx_z_1; // @[Bundles.scala 39:15]
  wire [20:0] tx_z_2 = tx_c + txInc_c; // @[Bundles.scala 38:17]
  wire [20:0] _tx_out_c_T_3 = |tx_z_2[20] ? 21'hfffff : tx_z_2; // @[Bundles.scala 39:15]
  wire [20:0] tx_z_3 = tx_d + txInc_d; // @[Bundles.scala 38:17]
  wire [20:0] _tx_out_d_T_3 = |tx_z_3[20] ? 21'hfffff : tx_z_3; // @[Bundles.scala 39:15]
  wire [20:0] tx_z_4 = tx_e + txInc_e; // @[Bundles.scala 38:17]
  wire [20:0] _tx_out_e_T_3 = |tx_z_4[20] ? 21'hfffff : tx_z_4; // @[Bundles.scala 39:15]
  wire [19:0] rxInc_a = {{19'd0}, _rxInc_a_T}; // @[RX.scala 87:19 RX.scala 89:9]
  wire [20:0] rx_z = rx_a + rxInc_a; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_a_T_3 = |rx_z[20] ? 21'hfffff : rx_z; // @[Bundles.scala 39:15]
  wire [19:0] rxInc_b = {{19'd0}, _rxInc_bT}; // @[RX.scala 87:19 RX.scala 89:9]
  wire [20:0] rx_z_1 = rx_b + rxInc_b; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_bT_3 = |rx_z_1[20] ? 21'hfffff : rx_z_1; // @[Bundles.scala 39:15]
  wire [19:0] rxInc_c = {{19'd0}, _rxInc_c_T}; // @[RX.scala 87:19 RX.scala 89:9]
  wire [20:0] rx_z_2 = rx_c + rxInc_c; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_c_T_3 = |rx_z_2[20] ? 21'hfffff : rx_z_2; // @[Bundles.scala 39:15]
  wire [19:0] rxInc_d = {{19'd0}, _rxInc_d_T}; // @[RX.scala 87:19 RX.scala 89:9]
  wire [20:0] rx_z_3 = rx_d + rxInc_d; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_d_T_3 = |rx_z_3[20] ? 21'hfffff : rx_z_3; // @[Bundles.scala 39:15]
  wire [19:0] rxInc_e = {{19'd0}, _rxInc_e_T}; // @[RX.scala 87:19 RX.scala 89:9]
  wire [20:0] rx_z_4 = rx_e + rxInc_e; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_e_T_3 = |rx_z_4[20] ? 21'hfffff : rx_z_4; // @[Bundles.scala 39:15]
  wire  txOut_ready = io_txc_source_io_enq_ready; // @[RX.scala 77:19 AsyncQueue.scala 217:19]
  wire [19:0] tx_out_1_a = _tx_out_a_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] tx_out_1_b = _tx_out_bT_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] tx_out_1_c = _tx_out_c_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] tx_out_1_d = _tx_out_d_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] tx_out_1_e = _tx_out_e_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire  rxOut_ready = io_rxc_source_io_enq_ready; // @[RX.scala 78:19 AsyncQueue.scala 217:19]
  wire [19:0] rx_out_1_a = _rx_out_a_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] rx_out_1_b = _rx_out_bT_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] rx_out_1_c = _rx_out_c_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] rx_out_1_d = _rx_out_d_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] rx_out_1_e = _rx_out_e_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  HellaQueue hqa ( // @[RX.scala 50:19]
    .clock(hqa_clock),
    .reset(hqa_reset),
    .io_enq_ready(hqa_io_enq_ready),
    .io_enq_valid(hqa_io_enq_valid),
    .io_enq_bits(hqa_io_enq_bits),
    .io_deq_ready(hqa_io_deq_ready),
    .io_deq_valid(hqa_io_deq_valid),
    .io_deq_bits(hqa_io_deq_bits)
  );
  HellaQueue hqb ( // @[RX.scala 51:19]
    .clock(hqb_clock),
    .reset(hqb_reset),
    .io_enq_ready(hqb_io_enq_ready),
    .io_enq_valid(hqb_io_enq_valid),
    .io_enq_bits(hqb_io_enq_bits),
    .io_deq_ready(hqb_io_deq_ready),
    .io_deq_valid(hqb_io_deq_valid),
    .io_deq_bits(hqb_io_deq_bits)
  );
  HellaQueue hqc ( // @[RX.scala 52:19]
    .clock(hqc_clock),
    .reset(hqc_reset),
    .io_enq_ready(hqc_io_enq_ready),
    .io_enq_valid(hqc_io_enq_valid),
    .io_enq_bits(hqc_io_enq_bits),
    .io_deq_ready(hqc_io_deq_ready),
    .io_deq_valid(hqc_io_deq_valid),
    .io_deq_bits(hqc_io_deq_bits)
  );
  HellaQueue hqd ( // @[RX.scala 53:19]
    .clock(hqd_clock),
    .reset(hqd_reset),
    .io_enq_ready(hqd_io_enq_ready),
    .io_enq_valid(hqd_io_enq_valid),
    .io_enq_bits(hqd_io_enq_bits),
    .io_deq_ready(hqd_io_deq_ready),
    .io_deq_valid(hqd_io_deq_valid),
    .io_deq_bits(hqd_io_deq_bits)
  );
  HellaQueue hqe ( // @[RX.scala 54:19]
    .clock(hqe_clock),
    .reset(hqe_reset),
    .io_enq_ready(hqe_io_enq_ready),
    .io_enq_valid(hqe_io_enq_valid),
    .io_enq_bits(hqe_io_enq_bits),
    .io_deq_ready(hqe_io_deq_ready),
    .io_deq_valid(hqe_io_deq_valid),
    .io_deq_bits(hqe_io_deq_bits)
  );
  AsyncQueueSource io_a_source ( // @[AsyncQueue.scala 216:24]
    .clock(io_a_source_clock),
    .reset(io_a_source_reset),
    .io_enq_ready(io_a_source_io_enq_ready),
    .io_enq_valid(io_a_source_io_enq_valid),
    .io_enq_bits(io_a_source_io_enq_bits),
    .io_async_mem_0(io_a_source_io_async_mem_0),
    .io_async_mem_1(io_a_source_io_async_mem_1),
    .io_async_mem_2(io_a_source_io_async_mem_2),
    .io_async_mem_3(io_a_source_io_async_mem_3),
    .io_async_mem_4(io_a_source_io_async_mem_4),
    .io_async_mem_5(io_a_source_io_async_mem_5),
    .io_async_mem_6(io_a_source_io_async_mem_6),
    .io_async_mem_7(io_a_source_io_async_mem_7),
    .io_async_ridx(io_a_source_io_async_ridx),
    .io_async_widx(io_a_source_io_async_widx),
    .io_async_safe_ridx_valid(io_a_source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(io_a_source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(io_a_source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(io_a_source_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource io_bsource ( // @[AsyncQueue.scala 216:24]
    .clock(io_bsource_clock),
    .reset(io_bsource_reset),
    .io_enq_ready(io_bsource_io_enq_ready),
    .io_enq_valid(io_bsource_io_enq_valid),
    .io_enq_bits(io_bsource_io_enq_bits),
    .io_async_mem_0(io_bsource_io_async_mem_0),
    .io_async_mem_1(io_bsource_io_async_mem_1),
    .io_async_mem_2(io_bsource_io_async_mem_2),
    .io_async_mem_3(io_bsource_io_async_mem_3),
    .io_async_mem_4(io_bsource_io_async_mem_4),
    .io_async_mem_5(io_bsource_io_async_mem_5),
    .io_async_mem_6(io_bsource_io_async_mem_6),
    .io_async_mem_7(io_bsource_io_async_mem_7),
    .io_async_ridx(io_bsource_io_async_ridx),
    .io_async_widx(io_bsource_io_async_widx),
    .io_async_safe_ridx_valid(io_bsource_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(io_bsource_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(io_bsource_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(io_bsource_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource io_c_source ( // @[AsyncQueue.scala 216:24]
    .clock(io_c_source_clock),
    .reset(io_c_source_reset),
    .io_enq_ready(io_c_source_io_enq_ready),
    .io_enq_valid(io_c_source_io_enq_valid),
    .io_enq_bits(io_c_source_io_enq_bits),
    .io_async_mem_0(io_c_source_io_async_mem_0),
    .io_async_mem_1(io_c_source_io_async_mem_1),
    .io_async_mem_2(io_c_source_io_async_mem_2),
    .io_async_mem_3(io_c_source_io_async_mem_3),
    .io_async_mem_4(io_c_source_io_async_mem_4),
    .io_async_mem_5(io_c_source_io_async_mem_5),
    .io_async_mem_6(io_c_source_io_async_mem_6),
    .io_async_mem_7(io_c_source_io_async_mem_7),
    .io_async_ridx(io_c_source_io_async_ridx),
    .io_async_widx(io_c_source_io_async_widx),
    .io_async_safe_ridx_valid(io_c_source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(io_c_source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(io_c_source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(io_c_source_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource io_d_source ( // @[AsyncQueue.scala 216:24]
    .clock(io_d_source_clock),
    .reset(io_d_source_reset),
    .io_enq_ready(io_d_source_io_enq_ready),
    .io_enq_valid(io_d_source_io_enq_valid),
    .io_enq_bits(io_d_source_io_enq_bits),
    .io_async_mem_0(io_d_source_io_async_mem_0),
    .io_async_mem_1(io_d_source_io_async_mem_1),
    .io_async_mem_2(io_d_source_io_async_mem_2),
    .io_async_mem_3(io_d_source_io_async_mem_3),
    .io_async_mem_4(io_d_source_io_async_mem_4),
    .io_async_mem_5(io_d_source_io_async_mem_5),
    .io_async_mem_6(io_d_source_io_async_mem_6),
    .io_async_mem_7(io_d_source_io_async_mem_7),
    .io_async_ridx(io_d_source_io_async_ridx),
    .io_async_widx(io_d_source_io_async_widx),
    .io_async_safe_ridx_valid(io_d_source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(io_d_source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(io_d_source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(io_d_source_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource io_e_source ( // @[AsyncQueue.scala 216:24]
    .clock(io_e_source_clock),
    .reset(io_e_source_reset),
    .io_enq_ready(io_e_source_io_enq_ready),
    .io_enq_valid(io_e_source_io_enq_valid),
    .io_enq_bits(io_e_source_io_enq_bits),
    .io_async_mem_0(io_e_source_io_async_mem_0),
    .io_async_mem_1(io_e_source_io_async_mem_1),
    .io_async_mem_2(io_e_source_io_async_mem_2),
    .io_async_mem_3(io_e_source_io_async_mem_3),
    .io_async_mem_4(io_e_source_io_async_mem_4),
    .io_async_mem_5(io_e_source_io_async_mem_5),
    .io_async_mem_6(io_e_source_io_async_mem_6),
    .io_async_mem_7(io_e_source_io_async_mem_7),
    .io_async_ridx(io_e_source_io_async_ridx),
    .io_async_widx(io_e_source_io_async_widx),
    .io_async_safe_ridx_valid(io_e_source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(io_e_source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(io_e_source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(io_e_source_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource_5 io_txc_source ( // @[AsyncQueue.scala 216:24]
    .clock(io_txc_source_clock),
    .reset(io_txc_source_reset),
    .io_enq_ready(io_txc_source_io_enq_ready),
    .io_enq_bits_a(io_txc_source_io_enq_bits_a),
    .io_enq_bits_b(io_txc_source_io_enq_bits_b),
    .io_enq_bits_c(io_txc_source_io_enq_bits_c),
    .io_enq_bits_d(io_txc_source_io_enq_bits_d),
    .io_enq_bits_e(io_txc_source_io_enq_bits_e),
    .io_async_mem_0_a(io_txc_source_io_async_mem_0_a),
    .io_async_mem_0_b(io_txc_source_io_async_mem_0_b),
    .io_async_mem_0_c(io_txc_source_io_async_mem_0_c),
    .io_async_mem_0_d(io_txc_source_io_async_mem_0_d),
    .io_async_mem_0_e(io_txc_source_io_async_mem_0_e),
    .io_async_ridx(io_txc_source_io_async_ridx),
    .io_async_widx(io_txc_source_io_async_widx),
    .io_async_safe_ridx_valid(io_txc_source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(io_txc_source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(io_txc_source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(io_txc_source_io_async_safe_sink_reset_n)
  );
  AsyncQueueSource_5 io_rxc_source ( // @[AsyncQueue.scala 216:24]
    .clock(io_rxc_source_clock),
    .reset(io_rxc_source_reset),
    .io_enq_ready(io_rxc_source_io_enq_ready),
    .io_enq_bits_a(io_rxc_source_io_enq_bits_a),
    .io_enq_bits_b(io_rxc_source_io_enq_bits_b),
    .io_enq_bits_c(io_rxc_source_io_enq_bits_c),
    .io_enq_bits_d(io_rxc_source_io_enq_bits_d),
    .io_enq_bits_e(io_rxc_source_io_enq_bits_e),
    .io_async_mem_0_a(io_rxc_source_io_async_mem_0_a),
    .io_async_mem_0_b(io_rxc_source_io_async_mem_0_b),
    .io_async_mem_0_c(io_rxc_source_io_async_mem_0_c),
    .io_async_mem_0_d(io_rxc_source_io_async_mem_0_d),
    .io_async_mem_0_e(io_rxc_source_io_async_mem_0_e),
    .io_async_ridx(io_rxc_source_io_async_ridx),
    .io_async_widx(io_rxc_source_io_async_widx),
    .io_async_safe_ridx_valid(io_rxc_source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(io_rxc_source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(io_rxc_source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(io_rxc_source_io_async_safe_sink_reset_n)
  );
  assign io_a_mem_0 = io_a_source_io_async_mem_0; // @[RX.scala 69:8]
  assign io_a_mem_1 = io_a_source_io_async_mem_1; // @[RX.scala 69:8]
  assign io_a_mem_2 = io_a_source_io_async_mem_2; // @[RX.scala 69:8]
  assign io_a_mem_3 = io_a_source_io_async_mem_3; // @[RX.scala 69:8]
  assign io_a_mem_4 = io_a_source_io_async_mem_4; // @[RX.scala 69:8]
  assign io_a_mem_5 = io_a_source_io_async_mem_5; // @[RX.scala 69:8]
  assign io_a_mem_6 = io_a_source_io_async_mem_6; // @[RX.scala 69:8]
  assign io_a_mem_7 = io_a_source_io_async_mem_7; // @[RX.scala 69:8]
  assign io_a_widx = io_a_source_io_async_widx; // @[RX.scala 69:8]
  assign io_a_safe_widx_valid = io_a_source_io_async_safe_widx_valid; // @[RX.scala 69:8]
  assign io_a_safe_source_reset_n = io_a_source_io_async_safe_source_reset_n; // @[RX.scala 69:8]
  assign io_bmem_0 = io_bsource_io_async_mem_0; // @[RX.scala 69:8]
  assign io_bmem_1 = io_bsource_io_async_mem_1; // @[RX.scala 69:8]
  assign io_bmem_2 = io_bsource_io_async_mem_2; // @[RX.scala 69:8]
  assign io_bmem_3 = io_bsource_io_async_mem_3; // @[RX.scala 69:8]
  assign io_bmem_4 = io_bsource_io_async_mem_4; // @[RX.scala 69:8]
  assign io_bmem_5 = io_bsource_io_async_mem_5; // @[RX.scala 69:8]
  assign io_bmem_6 = io_bsource_io_async_mem_6; // @[RX.scala 69:8]
  assign io_bmem_7 = io_bsource_io_async_mem_7; // @[RX.scala 69:8]
  assign io_bwidx = io_bsource_io_async_widx; // @[RX.scala 69:8]
  assign io_bsafe_widx_valid = io_bsource_io_async_safe_widx_valid; // @[RX.scala 69:8]
  assign io_bsafe_source_reset_n = io_bsource_io_async_safe_source_reset_n; // @[RX.scala 69:8]
  assign io_c_mem_0 = io_c_source_io_async_mem_0; // @[RX.scala 69:8]
  assign io_c_mem_1 = io_c_source_io_async_mem_1; // @[RX.scala 69:8]
  assign io_c_mem_2 = io_c_source_io_async_mem_2; // @[RX.scala 69:8]
  assign io_c_mem_3 = io_c_source_io_async_mem_3; // @[RX.scala 69:8]
  assign io_c_mem_4 = io_c_source_io_async_mem_4; // @[RX.scala 69:8]
  assign io_c_mem_5 = io_c_source_io_async_mem_5; // @[RX.scala 69:8]
  assign io_c_mem_6 = io_c_source_io_async_mem_6; // @[RX.scala 69:8]
  assign io_c_mem_7 = io_c_source_io_async_mem_7; // @[RX.scala 69:8]
  assign io_c_widx = io_c_source_io_async_widx; // @[RX.scala 69:8]
  assign io_c_safe_widx_valid = io_c_source_io_async_safe_widx_valid; // @[RX.scala 69:8]
  assign io_c_safe_source_reset_n = io_c_source_io_async_safe_source_reset_n; // @[RX.scala 69:8]
  assign io_d_mem_0 = io_d_source_io_async_mem_0; // @[RX.scala 69:8]
  assign io_d_mem_1 = io_d_source_io_async_mem_1; // @[RX.scala 69:8]
  assign io_d_mem_2 = io_d_source_io_async_mem_2; // @[RX.scala 69:8]
  assign io_d_mem_3 = io_d_source_io_async_mem_3; // @[RX.scala 69:8]
  assign io_d_mem_4 = io_d_source_io_async_mem_4; // @[RX.scala 69:8]
  assign io_d_mem_5 = io_d_source_io_async_mem_5; // @[RX.scala 69:8]
  assign io_d_mem_6 = io_d_source_io_async_mem_6; // @[RX.scala 69:8]
  assign io_d_mem_7 = io_d_source_io_async_mem_7; // @[RX.scala 69:8]
  assign io_d_widx = io_d_source_io_async_widx; // @[RX.scala 69:8]
  assign io_d_safe_widx_valid = io_d_source_io_async_safe_widx_valid; // @[RX.scala 69:8]
  assign io_d_safe_source_reset_n = io_d_source_io_async_safe_source_reset_n; // @[RX.scala 69:8]
  assign io_e_mem_0 = io_e_source_io_async_mem_0; // @[RX.scala 69:8]
  assign io_e_mem_1 = io_e_source_io_async_mem_1; // @[RX.scala 69:8]
  assign io_e_mem_2 = io_e_source_io_async_mem_2; // @[RX.scala 69:8]
  assign io_e_mem_3 = io_e_source_io_async_mem_3; // @[RX.scala 69:8]
  assign io_e_mem_4 = io_e_source_io_async_mem_4; // @[RX.scala 69:8]
  assign io_e_mem_5 = io_e_source_io_async_mem_5; // @[RX.scala 69:8]
  assign io_e_mem_6 = io_e_source_io_async_mem_6; // @[RX.scala 69:8]
  assign io_e_mem_7 = io_e_source_io_async_mem_7; // @[RX.scala 69:8]
  assign io_e_widx = io_e_source_io_async_widx; // @[RX.scala 69:8]
  assign io_e_safe_widx_valid = io_e_source_io_async_safe_widx_valid; // @[RX.scala 69:8]
  assign io_e_safe_source_reset_n = io_e_source_io_async_safe_source_reset_n; // @[RX.scala 69:8]
  assign io_rxc_mem_0_a = io_rxc_source_io_async_mem_0_a; // @[RX.scala 84:10]
  assign io_rxc_mem_0_b = io_rxc_source_io_async_mem_0_b; // @[RX.scala 84:10]
  assign io_rxc_mem_0_c = io_rxc_source_io_async_mem_0_c; // @[RX.scala 84:10]
  assign io_rxc_mem_0_d = io_rxc_source_io_async_mem_0_d; // @[RX.scala 84:10]
  assign io_rxc_mem_0_e = io_rxc_source_io_async_mem_0_e; // @[RX.scala 84:10]
  assign io_rxc_widx = io_rxc_source_io_async_widx; // @[RX.scala 84:10]
  assign io_rxc_safe_widx_valid = io_rxc_source_io_async_safe_widx_valid; // @[RX.scala 84:10]
  assign io_rxc_safe_source_reset_n = io_rxc_source_io_async_safe_source_reset_n; // @[RX.scala 84:10]
  assign io_txc_mem_0_a = io_txc_source_io_async_mem_0_a; // @[RX.scala 83:10]
  assign io_txc_mem_0_b = io_txc_source_io_async_mem_0_b; // @[RX.scala 83:10]
  assign io_txc_mem_0_c = io_txc_source_io_async_mem_0_c; // @[RX.scala 83:10]
  assign io_txc_mem_0_d = io_txc_source_io_async_mem_0_d; // @[RX.scala 83:10]
  assign io_txc_mem_0_e = io_txc_source_io_async_mem_0_e; // @[RX.scala 83:10]
  assign io_txc_widx = io_txc_source_io_async_widx; // @[RX.scala 83:10]
  assign io_txc_safe_widx_valid = io_txc_source_io_async_safe_widx_valid; // @[RX.scala 83:10]
  assign io_txc_safe_source_reset_n = io_txc_source_io_async_safe_source_reset_n; // @[RX.scala 83:10]
  assign hqa_clock = clock;
  assign hqa_reset = reset;
  assign hqa_io_enq_valid = b2c_data_valid & formatOH[0]; // @[RX.scala 62:35]
  assign hqa_io_enq_bits = b2c_data_concat; // @[RX.scala 37:18 RX.scala 38:14]
  assign hqa_io_deq_ready = io_a_source_io_enq_ready; // @[AsyncQueue.scala 217:19]
  assign hqb_clock = clock;
  assign hqb_reset = reset;
  assign hqb_io_enq_valid = b2c_data_valid & formatOH[1]; // @[RX.scala 62:35]
  assign hqb_io_enq_bits = b2c_data_concat; // @[RX.scala 37:18 RX.scala 38:14]
  assign hqb_io_deq_ready = io_bsource_io_enq_ready; // @[AsyncQueue.scala 217:19]
  assign hqc_clock = clock;
  assign hqc_reset = reset;
  assign hqc_io_enq_valid = b2c_data_valid & formatOH[2]; // @[RX.scala 62:35]
  assign hqc_io_enq_bits = b2c_data_concat; // @[RX.scala 37:18 RX.scala 38:14]
  assign hqc_io_deq_ready = io_c_source_io_enq_ready; // @[AsyncQueue.scala 217:19]
  assign hqd_clock = clock;
  assign hqd_reset = reset;
  assign hqd_io_enq_valid = b2c_data_valid & formatOH[3]; // @[RX.scala 62:35]
  assign hqd_io_enq_bits = b2c_data_concat; // @[RX.scala 37:18 RX.scala 38:14]
  assign hqd_io_deq_ready = io_d_source_io_enq_ready; // @[AsyncQueue.scala 217:19]
  assign hqe_clock = clock;
  assign hqe_reset = reset;
  assign hqe_io_enq_valid = b2c_data_valid & formatOH[4]; // @[RX.scala 62:35]
  assign hqe_io_enq_bits = b2c_data_concat; // @[RX.scala 37:18 RX.scala 38:14]
  assign hqe_io_deq_ready = io_e_source_io_enq_ready; // @[AsyncQueue.scala 217:19]
  assign io_a_source_clock = clock;
  assign io_a_source_reset = reset;
  assign io_a_source_io_enq_valid = hqa_io_deq_valid; // @[AsyncQueue.scala 217:19]
  assign io_a_source_io_enq_bits = hqa_io_deq_bits; // @[AsyncQueue.scala 217:19]
  assign io_a_source_io_async_ridx = io_a_ridx; // @[RX.scala 69:8]
  assign io_a_source_io_async_safe_ridx_valid = io_a_safe_ridx_valid; // @[RX.scala 69:8]
  assign io_a_source_io_async_safe_sink_reset_n = io_a_safe_sink_reset_n; // @[RX.scala 69:8]
  assign io_bsource_clock = clock;
  assign io_bsource_reset = reset;
  assign io_bsource_io_enq_valid = hqb_io_deq_valid; // @[AsyncQueue.scala 217:19]
  assign io_bsource_io_enq_bits = hqb_io_deq_bits; // @[AsyncQueue.scala 217:19]
  assign io_bsource_io_async_ridx = io_bridx; // @[RX.scala 69:8]
  assign io_bsource_io_async_safe_ridx_valid = io_bsafe_ridx_valid; // @[RX.scala 69:8]
  assign io_bsource_io_async_safe_sink_reset_n = io_bsafe_sink_reset_n; // @[RX.scala 69:8]
  assign io_c_source_clock = clock;
  assign io_c_source_reset = reset;
  assign io_c_source_io_enq_valid = hqc_io_deq_valid; // @[AsyncQueue.scala 217:19]
  assign io_c_source_io_enq_bits = hqc_io_deq_bits; // @[AsyncQueue.scala 217:19]
  assign io_c_source_io_async_ridx = io_c_ridx; // @[RX.scala 69:8]
  assign io_c_source_io_async_safe_ridx_valid = io_c_safe_ridx_valid; // @[RX.scala 69:8]
  assign io_c_source_io_async_safe_sink_reset_n = io_c_safe_sink_reset_n; // @[RX.scala 69:8]
  assign io_d_source_clock = clock;
  assign io_d_source_reset = reset;
  assign io_d_source_io_enq_valid = hqd_io_deq_valid; // @[AsyncQueue.scala 217:19]
  assign io_d_source_io_enq_bits = hqd_io_deq_bits; // @[AsyncQueue.scala 217:19]
  assign io_d_source_io_async_ridx = io_d_ridx; // @[RX.scala 69:8]
  assign io_d_source_io_async_safe_ridx_valid = io_d_safe_ridx_valid; // @[RX.scala 69:8]
  assign io_d_source_io_async_safe_sink_reset_n = io_d_safe_sink_reset_n; // @[RX.scala 69:8]
  assign io_e_source_clock = clock;
  assign io_e_source_reset = reset;
  assign io_e_source_io_enq_valid = hqe_io_deq_valid; // @[AsyncQueue.scala 217:19]
  assign io_e_source_io_enq_bits = hqe_io_deq_bits; // @[AsyncQueue.scala 217:19]
  assign io_e_source_io_async_ridx = io_e_ridx; // @[RX.scala 69:8]
  assign io_e_source_io_async_safe_ridx_valid = io_e_safe_ridx_valid; // @[RX.scala 69:8]
  assign io_e_source_io_async_safe_sink_reset_n = io_e_safe_sink_reset_n; // @[RX.scala 69:8]
  assign io_txc_source_clock = clock;
  assign io_txc_source_reset = reset;
  assign io_txc_source_io_enq_bits_a = tx_a; // @[RX.scala 77:19 RX.scala 81:14]
  assign io_txc_source_io_enq_bits_b = tx_b; // @[RX.scala 77:19 RX.scala 81:14]
  assign io_txc_source_io_enq_bits_c = tx_c; // @[RX.scala 77:19 RX.scala 81:14]
  assign io_txc_source_io_enq_bits_d = tx_d; // @[RX.scala 77:19 RX.scala 81:14]
  assign io_txc_source_io_enq_bits_e = tx_e; // @[RX.scala 77:19 RX.scala 81:14]
  assign io_txc_source_io_async_ridx = io_txc_ridx; // @[RX.scala 83:10]
  assign io_txc_source_io_async_safe_ridx_valid = io_txc_safe_ridx_valid; // @[RX.scala 83:10]
  assign io_txc_source_io_async_safe_sink_reset_n = io_txc_safe_sink_reset_n; // @[RX.scala 83:10]
  assign io_rxc_source_clock = clock;
  assign io_rxc_source_reset = reset;
  assign io_rxc_source_io_enq_bits_a = rx_a; // @[RX.scala 78:19 RX.scala 82:14]
  assign io_rxc_source_io_enq_bits_b = rx_b; // @[RX.scala 78:19 RX.scala 82:14]
  assign io_rxc_source_io_enq_bits_c = rx_c; // @[RX.scala 78:19 RX.scala 82:14]
  assign io_rxc_source_io_enq_bits_d = rx_d; // @[RX.scala 78:19 RX.scala 82:14]
  assign io_rxc_source_io_enq_bits_e = rx_e; // @[RX.scala 78:19 RX.scala 82:14]
  assign io_rxc_source_io_async_ridx = io_rxc_ridx; // @[RX.scala 84:10]
  assign io_rxc_source_io_async_safe_ridx_valid = io_rxc_safe_ridx_valid; // @[RX.scala 84:10]
  assign io_rxc_source_io_async_safe_sink_reset_n = io_rxc_safe_sink_reset_n; // @[RX.scala 84:10]
  always @(posedge clock) begin
    b2c_data_REG <= io_b2c_data; // @[RX.scala 24:33]
    b2c_data <= b2c_data_REG; // @[RX.scala 24:25]
    b2c_send_REG <= io_b2c_send; // @[RX.scala 25:33]
    if (reset) begin // @[RX.scala 25:25]
      b2c_send <= 1'h0; // @[RX.scala 25:25]
    end else begin
      b2c_send <= b2c_send_REG; // @[RX.scala 25:25]
    end
    if (reset) begin // @[RX.scala 27:24]
      beatCnt <= 2'h0; // @[RX.scala 27:24]
    end else if (b2c_send) begin // @[RX.scala 30:18]
      beatCnt <= _beatCnt_T_1; // @[RX.scala 31:13]
    end
    if (reset) begin // @[RX.scala 28:32]
      b2c_data_concat <= 32'h0; // @[RX.scala 28:32]
    end else begin
      b2c_data_concat <= _GEN_1[31:0];
    end
    if (reset) begin // @[RX.scala 29:31]
      b2c_data_valid <= 1'h0; // @[RX.scala 29:31]
    end else begin
      b2c_data_valid <= beatCnt == 2'h3; // @[RX.scala 34:18]
    end
    if (reset) begin // @[Parameters.scala 126:24]
      first_count <= 5'h0; // @[Parameters.scala 126:24]
    end else if (b2c_data_valid) begin // @[Parameters.scala 130:21]
      if (first) begin // @[Parameters.scala 130:35]
        if (3'h5 == first_beats_format) begin // @[Parameters.scala 129:54]
          first_count <= 5'h0; // @[Parameters.scala 129:54]
        end else begin
          first_count <= _GEN_6;
        end
      end else begin
        first_count <= _first_count_T_1;
      end
    end
    if (formatValid) begin // @[Reg.scala 16:19]
      format_r <= first_beats_format; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[RX.scala 73:19]
      tx_a <= 20'h0; // @[RX.scala 73:19]
    end else if (txOut_ready) begin // @[RX.scala 98:23]
      if (b2c_data_valid & formatOH[5]) begin // @[RX.scala 93:18]
        if (txInc_out_a_shiftAmount > 5'h14) begin // @[Bundles.scala 83:10]
          tx_a <= 20'hfffff;
        end else begin
          tx_a <= _txInc_out_a_T_3[20:1];
        end
      end else begin
        tx_a <= 20'h0;
      end
    end else begin
      tx_a <= tx_out_1_a; // @[RX.scala 96:6]
    end
    if (reset) begin // @[RX.scala 73:19]
      tx_b <= 20'h0; // @[RX.scala 73:19]
    end else if (txOut_ready) begin // @[RX.scala 98:23]
      if (b2c_data_valid & formatOH[5]) begin // @[RX.scala 93:18]
        if (txInc_out_bshiftAmount > 5'h14) begin // @[Bundles.scala 83:10]
          tx_b <= 20'hfffff;
        end else begin
          tx_b <= _txInc_out_bT_3[20:1];
        end
      end else begin
        tx_b <= 20'h0;
      end
    end else begin
      tx_b <= tx_out_1_b; // @[RX.scala 96:6]
    end
    if (reset) begin // @[RX.scala 73:19]
      tx_c <= 20'h0; // @[RX.scala 73:19]
    end else if (txOut_ready) begin // @[RX.scala 98:23]
      if (b2c_data_valid & formatOH[5]) begin // @[RX.scala 93:18]
        if (txInc_out_c_shiftAmount > 5'h14) begin // @[Bundles.scala 83:10]
          tx_c <= 20'hfffff;
        end else begin
          tx_c <= _txInc_out_c_T_3[20:1];
        end
      end else begin
        tx_c <= 20'h0;
      end
    end else begin
      tx_c <= tx_out_1_c; // @[RX.scala 96:6]
    end
    if (reset) begin // @[RX.scala 73:19]
      tx_d <= 20'h0; // @[RX.scala 73:19]
    end else if (txOut_ready) begin // @[RX.scala 98:23]
      if (b2c_data_valid & formatOH[5]) begin // @[RX.scala 93:18]
        if (txInc_out_d_shiftAmount > 5'h14) begin // @[Bundles.scala 83:10]
          tx_d <= 20'hfffff;
        end else begin
          tx_d <= _txInc_out_d_T_3[20:1];
        end
      end else begin
        tx_d <= 20'h0;
      end
    end else begin
      tx_d <= tx_out_1_d; // @[RX.scala 96:6]
    end
    if (reset) begin // @[RX.scala 73:19]
      tx_e <= 20'h0; // @[RX.scala 73:19]
    end else if (txOut_ready) begin // @[RX.scala 98:23]
      if (b2c_data_valid & formatOH[5]) begin // @[RX.scala 93:18]
        if (txInc_out_e_shiftAmount > 5'h14) begin // @[Bundles.scala 83:10]
          tx_e <= 20'hfffff;
        end else begin
          tx_e <= _txInc_out_e_T_3[20:1];
        end
      end else begin
        tx_e <= 20'h0;
      end
    end else begin
      tx_e <= tx_out_1_e; // @[RX.scala 96:6]
    end
    if (reset) begin // @[RX.scala 74:19]
      rx_a <= 20'h20; // @[RX.scala 74:19]
    end else if (rxOut_ready) begin // @[RX.scala 99:23]
      rx_a <= rxInc_a; // @[RX.scala 99:28]
    end else begin
      rx_a <= rx_out_1_a; // @[RX.scala 97:6]
    end
    if (reset) begin // @[RX.scala 74:19]
      rx_b <= 20'h20; // @[RX.scala 74:19]
    end else if (rxOut_ready) begin // @[RX.scala 99:23]
      rx_b <= rxInc_b; // @[RX.scala 99:28]
    end else begin
      rx_b <= rx_out_1_b; // @[RX.scala 97:6]
    end
    if (reset) begin // @[RX.scala 74:19]
      rx_c <= 20'h20; // @[RX.scala 74:19]
    end else if (rxOut_ready) begin // @[RX.scala 99:23]
      rx_c <= rxInc_c; // @[RX.scala 99:28]
    end else begin
      rx_c <= rx_out_1_c; // @[RX.scala 97:6]
    end
    if (reset) begin // @[RX.scala 74:19]
      rx_d <= 20'h20; // @[RX.scala 74:19]
    end else if (rxOut_ready) begin // @[RX.scala 99:23]
      rx_d <= rxInc_d; // @[RX.scala 99:28]
    end else begin
      rx_d <= rx_out_1_d; // @[RX.scala 97:6]
    end
    if (reset) begin // @[RX.scala 74:19]
      rx_e <= 20'h20; // @[RX.scala 74:19]
    end else if (rxOut_ready) begin // @[RX.scala 99:23]
      rx_e <= rxInc_e; // @[RX.scala 99:28]
    end else begin
      rx_e <= rx_out_1_e; // @[RX.scala 97:6]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~hqa_io_enq_valid | hqa_io_enq_ready | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at RX.scala:64 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"
            ); // @[RX.scala 64:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~hqa_io_enq_valid | hqa_io_enq_ready | reset)) begin
          $fatal; // @[RX.scala 64:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~hqb_io_enq_valid | hqb_io_enq_ready | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at RX.scala:64 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"
            ); // @[RX.scala 64:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~hqb_io_enq_valid | hqb_io_enq_ready | reset)) begin
          $fatal; // @[RX.scala 64:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~hqc_io_enq_valid | hqc_io_enq_ready | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at RX.scala:64 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"
            ); // @[RX.scala 64:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~hqc_io_enq_valid | hqc_io_enq_ready | reset)) begin
          $fatal; // @[RX.scala 64:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~hqd_io_enq_valid | hqd_io_enq_ready | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at RX.scala:64 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"
            ); // @[RX.scala 64:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~hqd_io_enq_valid | hqd_io_enq_ready | reset)) begin
          $fatal; // @[RX.scala 64:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~hqe_io_enq_valid | hqe_io_enq_ready | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at RX.scala:64 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"
            ); // @[RX.scala 64:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~hqe_io_enq_valid | hqe_io_enq_ready | reset)) begin
          $fatal; // @[RX.scala 64:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  b2c_data_REG = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  b2c_data = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  b2c_send_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  b2c_send = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  beatCnt = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  b2c_data_concat = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  b2c_data_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  first_count = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  format_r = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  tx_a = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  tx_b = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  tx_c = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  tx_d = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  tx_e = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  rx_a = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  rx_b = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  rx_c = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  rx_d = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  rx_e = _RAND_18[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncResetReg(
  output  io_q,
  input   io_clk,
  input   io_rst
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  reg_; // @[AsyncResetReg.scala 46:67]
  assign io_q = reg_; // @[AsyncResetReg.scala 50:8]
  always @(posedge io_clk or posedge io_rst) begin
    if (io_rst) begin
      reg_ <= 1'h1;
    end else begin
      reg_ <= 1'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  if (io_rst) begin
    reg_ = 1'h1;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockCrossingReg_w32(
  input         clock,
  input  [31:0] io_d,
  output [31:0] io_q,
  input         io_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cdc_reg; // @[Reg.scala 15:16]
  assign io_q = cdc_reg; // @[SynchronizerReg.scala 202:8]
  always @(posedge clock) begin
    if (io_en) begin // @[Reg.scala 16:19]
      cdc_reg <= io_d; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cdc_reg = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncQueueSink(
  input         clock,
  input         reset,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits,
  input  [31:0] io_async_mem_0,
  input  [31:0] io_async_mem_1,
  input  [31:0] io_async_mem_2,
  input  [31:0] io_async_mem_3,
  input  [31:0] io_async_mem_4,
  input  [31:0] io_async_mem_5,
  input  [31:0] io_async_mem_6,
  input  [31:0] io_async_mem_7,
  output [3:0]  io_async_ridx,
  input  [3:0]  io_async_widx,
  output        io_async_safe_ridx_valid,
  input         io_async_safe_widx_valid,
  input         io_async_safe_source_reset_n,
  output        io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  widx_widx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  widx_widx_gray_reset; // @[ShiftReg.scala 45:23]
  wire [3:0] widx_widx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire [3:0] widx_widx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  io_deq_bits_deq_bits_reg_clock; // @[SynchronizerReg.scala 207:25]
  wire [31:0] io_deq_bits_deq_bits_reg_io_d; // @[SynchronizerReg.scala 207:25]
  wire [31:0] io_deq_bits_deq_bits_reg_io_q; // @[SynchronizerReg.scala 207:25]
  wire  io_deq_bits_deq_bits_reg_io_en; // @[SynchronizerReg.scala 207:25]
  wire  sink_valid_0_io_in; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_io_out; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_clock; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_reset; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_1_io_in; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_io_out; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_clock; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_reset; // @[AsyncQueue.scala 169:33]
  wire  source_extend_io_in; // @[AsyncQueue.scala 171:31]
  wire  source_extend_io_out; // @[AsyncQueue.scala 171:31]
  wire  source_extend_clock; // @[AsyncQueue.scala 171:31]
  wire  source_extend_reset; // @[AsyncQueue.scala 171:31]
  wire  source_valid_io_in; // @[AsyncQueue.scala 172:31]
  wire  source_valid_io_out; // @[AsyncQueue.scala 172:31]
  wire  source_valid_clock; // @[AsyncQueue.scala 172:31]
  wire  source_valid_reset; // @[AsyncQueue.scala 172:31]
  wire  _ridx_T_1 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  source_ready = source_valid_io_out;
  wire  _ridx_T_2 = ~source_ready; // @[AsyncQueue.scala 144:79]
  reg [3:0] ridx_ridx_bin; // @[AsyncQueue.scala 52:25]
  wire [3:0] _GEN_8 = {{3'd0}, _ridx_T_1}; // @[AsyncQueue.scala 53:43]
  wire [3:0] _ridx_incremented_T_1 = ridx_ridx_bin + _GEN_8; // @[AsyncQueue.scala 53:43]
  wire [3:0] ridx_incremented = _ridx_T_2 ? 4'h0 : _ridx_incremented_T_1; // @[AsyncQueue.scala 53:23]
  wire [3:0] _GEN_9 = {{1'd0}, ridx_incremented[3:1]}; // @[AsyncQueue.scala 54:17]
  wire [3:0] ridx = ridx_incremented ^ _GEN_9; // @[AsyncQueue.scala 54:17]
  wire [3:0] widx = widx_widx_gray_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire [2:0] _index_T_2 = {ridx[3], 2'h0}; // @[AsyncQueue.scala 152:75]
  wire [2:0] index = ridx[2:0] ^ _index_T_2; // @[AsyncQueue.scala 152:55]
  wire [31:0] _GEN_1 = 3'h1 == index ? io_async_mem_1 : io_async_mem_0; // @[SynchronizerReg.scala 209:18 SynchronizerReg.scala 209:18]
  wire [31:0] _GEN_2 = 3'h2 == index ? io_async_mem_2 : _GEN_1; // @[SynchronizerReg.scala 209:18 SynchronizerReg.scala 209:18]
  wire [31:0] _GEN_3 = 3'h3 == index ? io_async_mem_3 : _GEN_2; // @[SynchronizerReg.scala 209:18 SynchronizerReg.scala 209:18]
  wire [31:0] _GEN_4 = 3'h4 == index ? io_async_mem_4 : _GEN_3; // @[SynchronizerReg.scala 209:18 SynchronizerReg.scala 209:18]
  wire [31:0] _GEN_5 = 3'h5 == index ? io_async_mem_5 : _GEN_4; // @[SynchronizerReg.scala 209:18 SynchronizerReg.scala 209:18]
  wire [31:0] _GEN_6 = 3'h6 == index ? io_async_mem_6 : _GEN_5; // @[SynchronizerReg.scala 209:18 SynchronizerReg.scala 209:18]
  reg  valid_reg; // @[AsyncQueue.scala 161:56]
  reg [3:0] ridx_gray; // @[AsyncQueue.scala 164:55]
  AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_widx_gray ( // @[ShiftReg.scala 45:23]
    .clock(widx_widx_gray_clock),
    .reset(widx_widx_gray_reset),
    .io_d(widx_widx_gray_io_d),
    .io_q(widx_widx_gray_io_q)
  );
  ClockCrossingReg_w32 io_deq_bits_deq_bits_reg ( // @[SynchronizerReg.scala 207:25]
    .clock(io_deq_bits_deq_bits_reg_clock),
    .io_d(io_deq_bits_deq_bits_reg_io_d),
    .io_q(io_deq_bits_deq_bits_reg_io_q),
    .io_en(io_deq_bits_deq_bits_reg_io_en)
  );
  AsyncValidSync sink_valid_0 ( // @[AsyncQueue.scala 168:33]
    .io_in(sink_valid_0_io_in),
    .io_out(sink_valid_0_io_out),
    .clock(sink_valid_0_clock),
    .reset(sink_valid_0_reset)
  );
  AsyncValidSync sink_valid_1 ( // @[AsyncQueue.scala 169:33]
    .io_in(sink_valid_1_io_in),
    .io_out(sink_valid_1_io_out),
    .clock(sink_valid_1_clock),
    .reset(sink_valid_1_reset)
  );
  AsyncValidSync source_extend ( // @[AsyncQueue.scala 171:31]
    .io_in(source_extend_io_in),
    .io_out(source_extend_io_out),
    .clock(source_extend_clock),
    .reset(source_extend_reset)
  );
  AsyncValidSync source_valid ( // @[AsyncQueue.scala 172:31]
    .io_in(source_valid_io_in),
    .io_out(source_valid_io_out),
    .clock(source_valid_clock),
    .reset(source_valid_reset)
  );
  assign io_deq_valid = valid_reg & source_ready; // @[AsyncQueue.scala 162:29]
  assign io_deq_bits = io_deq_bits_deq_bits_reg_io_q; // @[SynchronizerReg.scala 211:26 SynchronizerReg.scala 211:26]
  assign io_async_ridx = ridx_gray; // @[AsyncQueue.scala 165:17]
  assign io_async_safe_ridx_valid = sink_valid_1_io_out; // @[AsyncQueue.scala 185:20]
  assign io_async_safe_sink_reset_n = ~reset; // @[AsyncQueue.scala 189:25]
  assign widx_widx_gray_clock = clock;
  assign widx_widx_gray_reset = reset;
  assign widx_widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 47:16]
  assign io_deq_bits_deq_bits_reg_clock = clock;
  assign io_deq_bits_deq_bits_reg_io_d = 3'h7 == index ? io_async_mem_7 : _GEN_6; // @[SynchronizerReg.scala 209:18 SynchronizerReg.scala 209:18]
  assign io_deq_bits_deq_bits_reg_io_en = source_ready & ridx != widx; // @[AsyncQueue.scala 146:28]
  assign sink_valid_0_io_in = 1'h1; // @[AsyncQueue.scala 183:24]
  assign sink_valid_0_clock = clock; // @[AsyncQueue.scala 178:25]
  assign sink_valid_0_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 173:66]
  assign sink_valid_1_io_in = sink_valid_0_io_out; // @[AsyncQueue.scala 184:24]
  assign sink_valid_1_clock = clock; // @[AsyncQueue.scala 179:25]
  assign sink_valid_1_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 174:66]
  assign source_extend_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 186:25]
  assign source_extend_clock = clock; // @[AsyncQueue.scala 180:25]
  assign source_extend_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 175:66]
  assign source_valid_io_in = source_extend_io_out; // @[AsyncQueue.scala 187:24]
  assign source_valid_clock = clock; // @[AsyncQueue.scala 181:25]
  assign source_valid_reset = reset; // @[AsyncQueue.scala 176:34]
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ridx_ridx_bin <= 4'h0;
    end else if (_ridx_T_2) begin
      ridx_ridx_bin <= 4'h0;
    end else begin
      ridx_ridx_bin <= _ridx_incremented_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      valid_reg <= 1'h0;
    end else begin
      valid_reg <= source_ready & ridx != widx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ridx_gray <= 4'h0;
    end else begin
      ridx_gray <= ridx_incremented ^ _GEN_9;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ridx_ridx_bin = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ridx_gray = _RAND_2[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ridx_ridx_bin = 4'h0;
  end
  if (reset) begin
    valid_reg = 1'h0;
  end
  if (reset) begin
    ridx_gray = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockCrossingReg_w100(
  input         clock,
  input  [99:0] io_d,
  output [99:0] io_q,
  input         io_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [99:0] cdc_reg; // @[Reg.scala 15:16]
  assign io_q = cdc_reg; // @[SynchronizerReg.scala 202:8]
  always @(posedge clock) begin
    if (io_en) begin // @[Reg.scala 16:19]
      cdc_reg <= io_d; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  cdc_reg = _RAND_0[99:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncQueueSink_5(
  input         clock,
  input         reset,
  input         io_deq_ready,
  output        io_deq_valid,
  output [19:0] io_deq_bits_a,
  output [19:0] io_deq_bits_b,
  output [19:0] io_deq_bits_c,
  output [19:0] io_deq_bits_d,
  output [19:0] io_deq_bits_e,
  input  [19:0] io_async_mem_0_a,
  input  [19:0] io_async_mem_0_b,
  input  [19:0] io_async_mem_0_c,
  input  [19:0] io_async_mem_0_d,
  input  [19:0] io_async_mem_0_e,
  output        io_async_ridx,
  input         io_async_widx,
  output        io_async_safe_ridx_valid,
  input         io_async_safe_widx_valid,
  input         io_async_safe_source_reset_n,
  output        io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  widx_widx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  widx_widx_gray_reset; // @[ShiftReg.scala 45:23]
  wire  widx_widx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire  widx_widx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  io_deq_bits_deq_bits_reg_clock; // @[SynchronizerReg.scala 207:25]
  wire [99:0] io_deq_bits_deq_bits_reg_io_d; // @[SynchronizerReg.scala 207:25]
  wire [99:0] io_deq_bits_deq_bits_reg_io_q; // @[SynchronizerReg.scala 207:25]
  wire  io_deq_bits_deq_bits_reg_io_en; // @[SynchronizerReg.scala 207:25]
  wire  sink_valid_0_io_in; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_io_out; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_clock; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_reset; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_1_io_in; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_io_out; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_clock; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_reset; // @[AsyncQueue.scala 169:33]
  wire  source_extend_io_in; // @[AsyncQueue.scala 171:31]
  wire  source_extend_io_out; // @[AsyncQueue.scala 171:31]
  wire  source_extend_clock; // @[AsyncQueue.scala 171:31]
  wire  source_extend_reset; // @[AsyncQueue.scala 171:31]
  wire  source_valid_io_in; // @[AsyncQueue.scala 172:31]
  wire  source_valid_io_out; // @[AsyncQueue.scala 172:31]
  wire  source_valid_clock; // @[AsyncQueue.scala 172:31]
  wire  source_valid_reset; // @[AsyncQueue.scala 172:31]
  wire  source_ready = source_valid_io_out;
  wire  _ridx_T_2 = ~source_ready; // @[AsyncQueue.scala 144:79]
  reg  ridx_ridx_bin; // @[AsyncQueue.scala 52:25]
  wire  ridx_incremented = _ridx_T_2 ? 1'h0 : ridx_ridx_bin + io_deq_valid; // @[AsyncQueue.scala 53:23]
  wire  widx = widx_widx_gray_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire [39:0] io_deq_bits_deq_bits_reg_io_d_lo = {io_async_mem_0_d,io_async_mem_0_e}; // @[SynchronizerReg.scala 209:24]
  wire [59:0] io_deq_bits_deq_bits_reg_io_d_hi = {io_async_mem_0_a,io_async_mem_0_b,io_async_mem_0_c}; // @[SynchronizerReg.scala 209:24]
  wire [99:0] _io_deq_bits_WIRE_1 = io_deq_bits_deq_bits_reg_io_q;
  reg  valid_reg; // @[AsyncQueue.scala 161:56]
  reg  ridx_gray; // @[AsyncQueue.scala 164:55]
  AsyncResetSynchronizerShiftReg_w1_d3_i0_20 widx_widx_gray ( // @[ShiftReg.scala 45:23]
    .clock(widx_widx_gray_clock),
    .reset(widx_widx_gray_reset),
    .io_d(widx_widx_gray_io_d),
    .io_q(widx_widx_gray_io_q)
  );
  ClockCrossingReg_w100 io_deq_bits_deq_bits_reg ( // @[SynchronizerReg.scala 207:25]
    .clock(io_deq_bits_deq_bits_reg_clock),
    .io_d(io_deq_bits_deq_bits_reg_io_d),
    .io_q(io_deq_bits_deq_bits_reg_io_q),
    .io_en(io_deq_bits_deq_bits_reg_io_en)
  );
  AsyncValidSync sink_valid_0 ( // @[AsyncQueue.scala 168:33]
    .io_in(sink_valid_0_io_in),
    .io_out(sink_valid_0_io_out),
    .clock(sink_valid_0_clock),
    .reset(sink_valid_0_reset)
  );
  AsyncValidSync sink_valid_1 ( // @[AsyncQueue.scala 169:33]
    .io_in(sink_valid_1_io_in),
    .io_out(sink_valid_1_io_out),
    .clock(sink_valid_1_clock),
    .reset(sink_valid_1_reset)
  );
  AsyncValidSync source_extend ( // @[AsyncQueue.scala 171:31]
    .io_in(source_extend_io_in),
    .io_out(source_extend_io_out),
    .clock(source_extend_clock),
    .reset(source_extend_reset)
  );
  AsyncValidSync source_valid ( // @[AsyncQueue.scala 172:31]
    .io_in(source_valid_io_in),
    .io_out(source_valid_io_out),
    .clock(source_valid_clock),
    .reset(source_valid_reset)
  );
  assign io_deq_valid = valid_reg & source_ready; // @[AsyncQueue.scala 162:29]
  assign io_deq_bits_a = _io_deq_bits_WIRE_1[99:80]; // @[SynchronizerReg.scala 211:26]
  assign io_deq_bits_b = _io_deq_bits_WIRE_1[79:60]; // @[SynchronizerReg.scala 211:26]
  assign io_deq_bits_c = _io_deq_bits_WIRE_1[59:40]; // @[SynchronizerReg.scala 211:26]
  assign io_deq_bits_d = _io_deq_bits_WIRE_1[39:20]; // @[SynchronizerReg.scala 211:26]
  assign io_deq_bits_e = _io_deq_bits_WIRE_1[19:0]; // @[SynchronizerReg.scala 211:26]
  assign io_async_ridx = ridx_gray; // @[AsyncQueue.scala 165:17]
  assign io_async_safe_ridx_valid = sink_valid_1_io_out; // @[AsyncQueue.scala 185:20]
  assign io_async_safe_sink_reset_n = ~reset; // @[AsyncQueue.scala 189:25]
  assign widx_widx_gray_clock = clock;
  assign widx_widx_gray_reset = reset;
  assign widx_widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 47:16]
  assign io_deq_bits_deq_bits_reg_clock = clock;
  assign io_deq_bits_deq_bits_reg_io_d = {io_deq_bits_deq_bits_reg_io_d_hi,io_deq_bits_deq_bits_reg_io_d_lo}; // @[SynchronizerReg.scala 209:24]
  assign io_deq_bits_deq_bits_reg_io_en = source_ready & ridx_incremented != widx; // @[AsyncQueue.scala 146:28]
  assign sink_valid_0_io_in = 1'h1; // @[AsyncQueue.scala 183:24]
  assign sink_valid_0_clock = clock; // @[AsyncQueue.scala 178:25]
  assign sink_valid_0_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 173:66]
  assign sink_valid_1_io_in = sink_valid_0_io_out; // @[AsyncQueue.scala 184:24]
  assign sink_valid_1_clock = clock; // @[AsyncQueue.scala 179:25]
  assign sink_valid_1_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 174:66]
  assign source_extend_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 186:25]
  assign source_extend_clock = clock; // @[AsyncQueue.scala 180:25]
  assign source_extend_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 175:66]
  assign source_valid_io_in = source_extend_io_out; // @[AsyncQueue.scala 187:24]
  assign source_valid_clock = clock; // @[AsyncQueue.scala 181:25]
  assign source_valid_reset = reset; // @[AsyncQueue.scala 176:34]
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ridx_ridx_bin <= 1'h0;
    end else if (_ridx_T_2) begin
      ridx_ridx_bin <= 1'h0;
    end else begin
      ridx_ridx_bin <= ridx_ridx_bin + io_deq_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      valid_reg <= 1'h0;
    end else begin
      valid_reg <= source_ready & ridx_incremented != widx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ridx_gray <= 1'h0;
    end else if (_ridx_T_2) begin
      ridx_gray <= 1'h0;
    end else begin
      ridx_gray <= ridx_ridx_bin + io_deq_valid;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ridx_ridx_bin = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ridx_gray = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ridx_ridx_bin = 1'h0;
  end
  if (reset) begin
    valid_reg = 1'h0;
  end
  if (reset) begin
    ridx_gray = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ShiftQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input  [6:0]  io_enq_bits_beats,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last,
  output [6:0]  io_deq_bits_beats
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  valid_0; // @[ShiftQueue.scala 21:30]
  reg  valid_1; // @[ShiftQueue.scala 21:30]
  reg [31:0] elts_0_data; // @[ShiftQueue.scala 22:25]
  reg  elts_0_last; // @[ShiftQueue.scala 22:25]
  reg [6:0] elts_0_beats; // @[ShiftQueue.scala 22:25]
  reg [31:0] elts_1_data; // @[ShiftQueue.scala 22:25]
  reg  elts_1_last; // @[ShiftQueue.scala 22:25]
  reg [6:0] elts_1_beats; // @[ShiftQueue.scala 22:25]
  wire  _wen_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _wen_T_3 = valid_1 | _wen_T; // @[ShiftQueue.scala 30:28]
  wire  _wen_T_7 = _wen_T & ~valid_0; // @[ShiftQueue.scala 31:45]
  wire  wen = io_deq_ready ? _wen_T_3 : _wen_T_7; // @[ShiftQueue.scala 29:10]
  wire  _valid_0_T_6 = _wen_T | valid_0; // @[ShiftQueue.scala 37:45]
  wire  _wen_T_10 = _wen_T & valid_1; // @[ShiftQueue.scala 30:45]
  wire  _wen_T_13 = _wen_T & valid_0; // @[ShiftQueue.scala 31:25]
  wire  _wen_T_15 = _wen_T & valid_0 & ~valid_1; // @[ShiftQueue.scala 31:45]
  wire  wen_1 = io_deq_ready ? _wen_T_10 : _wen_T_15; // @[ShiftQueue.scala 29:10]
  wire  _valid_1_T_6 = _wen_T_13 | valid_1; // @[ShiftQueue.scala 37:45]
  assign io_enq_ready = ~valid_1; // @[ShiftQueue.scala 40:19]
  assign io_deq_valid = valid_0; // @[ShiftQueue.scala 41:16]
  assign io_deq_bits_data = elts_0_data; // @[ShiftQueue.scala 42:15]
  assign io_deq_bits_last = elts_0_last; // @[ShiftQueue.scala 42:15]
  assign io_deq_bits_beats = elts_0_beats; // @[ShiftQueue.scala 42:15]
  always @(posedge clock) begin
    if (reset) begin // @[ShiftQueue.scala 21:30]
      valid_0 <= 1'h0; // @[ShiftQueue.scala 21:30]
    end else if (io_deq_ready) begin // @[ShiftQueue.scala 35:10]
      valid_0 <= _wen_T_3;
    end else begin
      valid_0 <= _valid_0_T_6;
    end
    if (reset) begin // @[ShiftQueue.scala 21:30]
      valid_1 <= 1'h0; // @[ShiftQueue.scala 21:30]
    end else if (io_deq_ready) begin // @[ShiftQueue.scala 35:10]
      valid_1 <= _wen_T_10;
    end else begin
      valid_1 <= _valid_1_T_6;
    end
    if (wen) begin // @[ShiftQueue.scala 32:16]
      if (valid_1) begin // @[ShiftQueue.scala 27:57]
        elts_0_data <= elts_1_data;
      end else begin
        elts_0_data <= io_enq_bits_data;
      end
    end
    if (wen) begin // @[ShiftQueue.scala 32:16]
      if (valid_1) begin // @[ShiftQueue.scala 27:57]
        elts_0_last <= elts_1_last;
      end else begin
        elts_0_last <= io_enq_bits_last;
      end
    end
    if (wen) begin // @[ShiftQueue.scala 32:16]
      if (valid_1) begin // @[ShiftQueue.scala 27:57]
        elts_0_beats <= elts_1_beats;
      end else begin
        elts_0_beats <= io_enq_bits_beats;
      end
    end
    if (wen_1) begin // @[ShiftQueue.scala 32:16]
      elts_1_data <= io_enq_bits_data; // @[ShiftQueue.scala 32:26]
    end
    if (wen_1) begin // @[ShiftQueue.scala 32:16]
      elts_1_last <= io_enq_bits_last; // @[ShiftQueue.scala 32:26]
    end
    if (wen_1) begin // @[ShiftQueue.scala 32:16]
      elts_1_beats <= io_enq_bits_beats; // @[ShiftQueue.scala 32:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  valid_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  elts_0_data = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  elts_0_last = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  elts_0_beats = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  elts_1_data = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  elts_1_last = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  elts_1_beats = _RAND_7[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TX(
  input         clock,
  input         reset,
  output        io_c2b_clk,
  output        io_c2b_rst,
  output        io_c2b_send,
  output [7:0]  io_c2b_data,
  output        io_sa_ready,
  input         io_sa_valid,
  input  [31:0] io_sa_bits_data,
  input         io_sa_bits_last,
  input  [6:0]  io_sa_bits_beats,
  output        io_sb_ready,
  input  [31:0] io_sb_bits_data,
  input         io_sb_bits_last,
  output        io_sc_ready,
  input  [31:0] io_sc_bits_data,
  input         io_sc_bits_last,
  output        io_sd_ready,
  input         io_sd_valid,
  input  [31:0] io_sd_bits_data,
  input         io_sd_bits_last,
  input  [6:0]  io_sd_bits_beats,
  input  [31:0] io_se_bits_data,
  input  [19:0] io_rxc_mem_0_a,
  input  [19:0] io_rxc_mem_0_b,
  input  [19:0] io_rxc_mem_0_c,
  input  [19:0] io_rxc_mem_0_d,
  input  [19:0] io_rxc_mem_0_e,
  output        io_rxc_ridx,
  input         io_rxc_widx,
  output        io_rxc_safe_ridx_valid,
  input         io_rxc_safe_widx_valid,
  input         io_rxc_safe_source_reset_n,
  output        io_rxc_safe_sink_reset_n,
  input  [19:0] io_txc_mem_0_a,
  input  [19:0] io_txc_mem_0_b,
  input  [19:0] io_txc_mem_0_c,
  input  [19:0] io_txc_mem_0_d,
  input  [19:0] io_txc_mem_0_e,
  output        io_txc_ridx,
  input         io_txc_widx,
  output        io_txc_safe_ridx_valid,
  input         io_txc_safe_widx_valid,
  input         io_txc_safe_source_reset_n,
  output        io_txc_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  wire  rxInc_sink_clock; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_reset; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_io_deq_ready; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_io_deq_valid; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_deq_bits_a; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_deq_bits_b; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_deq_bits_c; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_deq_bits_d; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_deq_bits_e; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_async_mem_0_a; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_async_mem_0_b; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_async_mem_0_c; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_async_mem_0_d; // @[AsyncQueue.scala 207:22]
  wire [19:0] rxInc_sink_io_async_mem_0_e; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_io_async_ridx; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_io_async_widx; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 207:22]
  wire  rxInc_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_clock; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_reset; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_io_deq_ready; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_io_deq_valid; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_deq_bits_a; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_deq_bits_b; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_deq_bits_c; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_deq_bits_d; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_deq_bits_e; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_async_mem_0_a; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_async_mem_0_b; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_async_mem_0_c; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_async_mem_0_d; // @[AsyncQueue.scala 207:22]
  wire [19:0] txInc_sink_io_async_mem_0_e; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_io_async_ridx; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_io_async_widx; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 207:22]
  wire  txInc_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 207:22]
  wire  qa_q_clock; // @[ShiftQueue.scala 60:19]
  wire  qa_q_reset; // @[ShiftQueue.scala 60:19]
  wire  qa_q_io_enq_ready; // @[ShiftQueue.scala 60:19]
  wire  qa_q_io_enq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qa_q_io_enq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qa_q_io_enq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qa_q_io_enq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qa_q_io_deq_ready; // @[ShiftQueue.scala 60:19]
  wire  qa_q_io_deq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qa_q_io_deq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qa_q_io_deq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qa_q_io_deq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qb_q_clock; // @[ShiftQueue.scala 60:19]
  wire  qb_q_reset; // @[ShiftQueue.scala 60:19]
  wire  qb_q_io_enq_ready; // @[ShiftQueue.scala 60:19]
  wire  qb_q_io_enq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qb_q_io_enq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qb_q_io_enq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qb_q_io_enq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qb_q_io_deq_ready; // @[ShiftQueue.scala 60:19]
  wire  qb_q_io_deq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qb_q_io_deq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qb_q_io_deq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qb_q_io_deq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qc_q_clock; // @[ShiftQueue.scala 60:19]
  wire  qc_q_reset; // @[ShiftQueue.scala 60:19]
  wire  qc_q_io_enq_ready; // @[ShiftQueue.scala 60:19]
  wire  qc_q_io_enq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qc_q_io_enq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qc_q_io_enq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qc_q_io_enq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qc_q_io_deq_ready; // @[ShiftQueue.scala 60:19]
  wire  qc_q_io_deq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qc_q_io_deq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qc_q_io_deq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qc_q_io_deq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qd_q_clock; // @[ShiftQueue.scala 60:19]
  wire  qd_q_reset; // @[ShiftQueue.scala 60:19]
  wire  qd_q_io_enq_ready; // @[ShiftQueue.scala 60:19]
  wire  qd_q_io_enq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qd_q_io_enq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qd_q_io_enq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qd_q_io_enq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qd_q_io_deq_ready; // @[ShiftQueue.scala 60:19]
  wire  qd_q_io_deq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qd_q_io_deq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qd_q_io_deq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qd_q_io_deq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qe_q_clock; // @[ShiftQueue.scala 60:19]
  wire  qe_q_reset; // @[ShiftQueue.scala 60:19]
  wire  qe_q_io_enq_ready; // @[ShiftQueue.scala 60:19]
  wire  qe_q_io_enq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qe_q_io_enq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qe_q_io_enq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qe_q_io_enq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  qe_q_io_deq_ready; // @[ShiftQueue.scala 60:19]
  wire  qe_q_io_deq_valid; // @[ShiftQueue.scala 60:19]
  wire [31:0] qe_q_io_deq_bits_data; // @[ShiftQueue.scala 60:19]
  wire  qe_q_io_deq_bits_last; // @[ShiftQueue.scala 60:19]
  wire [6:0] qe_q_io_deq_bits_beats; // @[ShiftQueue.scala 60:19]
  wire  ioX_cq_clock; // @[TX.scala 56:20]
  wire  ioX_cq_reset; // @[TX.scala 56:20]
  wire  ioX_cq_io_enq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_io_enq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_io_enq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_io_enq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_io_enq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_io_deq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_io_deq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_io_deq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_io_deq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_io_deq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_1_clock; // @[TX.scala 56:20]
  wire  ioX_cq_1_reset; // @[TX.scala 56:20]
  wire  ioX_cq_1_io_enq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_1_io_enq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_1_io_enq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_1_io_enq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_1_io_enq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_1_io_deq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_1_io_deq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_1_io_deq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_1_io_deq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_1_io_deq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_2_clock; // @[TX.scala 56:20]
  wire  ioX_cq_2_reset; // @[TX.scala 56:20]
  wire  ioX_cq_2_io_enq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_2_io_enq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_2_io_enq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_2_io_enq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_2_io_enq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_2_io_deq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_2_io_deq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_2_io_deq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_2_io_deq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_2_io_deq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_3_clock; // @[TX.scala 56:20]
  wire  ioX_cq_3_reset; // @[TX.scala 56:20]
  wire  ioX_cq_3_io_enq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_3_io_enq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_3_io_enq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_3_io_enq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_3_io_enq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_3_io_deq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_3_io_deq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_3_io_deq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_3_io_deq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_3_io_deq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_4_clock; // @[TX.scala 56:20]
  wire  ioX_cq_4_reset; // @[TX.scala 56:20]
  wire  ioX_cq_4_io_enq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_4_io_enq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_4_io_enq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_4_io_enq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_4_io_enq_bits_beats; // @[TX.scala 56:20]
  wire  ioX_cq_4_io_deq_ready; // @[TX.scala 56:20]
  wire  ioX_cq_4_io_deq_valid; // @[TX.scala 56:20]
  wire [31:0] ioX_cq_4_io_deq_bits_data; // @[TX.scala 56:20]
  wire  ioX_cq_4_io_deq_bits_last; // @[TX.scala 56:20]
  wire [6:0] ioX_cq_4_io_deq_bits_beats; // @[TX.scala 56:20]
  wire  rxQ_clock; // @[TX.scala 64:19]
  wire  rxQ_reset; // @[TX.scala 64:19]
  wire  rxQ_io_enq_ready; // @[TX.scala 64:19]
  wire  rxQ_io_enq_valid; // @[TX.scala 64:19]
  wire [31:0] rxQ_io_enq_bits_data; // @[TX.scala 64:19]
  wire  rxQ_io_enq_bits_last; // @[TX.scala 64:19]
  wire [6:0] rxQ_io_enq_bits_beats; // @[TX.scala 64:19]
  wire  rxQ_io_deq_ready; // @[TX.scala 64:19]
  wire  rxQ_io_deq_valid; // @[TX.scala 64:19]
  wire [31:0] rxQ_io_deq_bits_data; // @[TX.scala 64:19]
  wire  rxQ_io_deq_bits_last; // @[TX.scala 64:19]
  wire [6:0] rxQ_io_deq_bits_beats; // @[TX.scala 64:19]
  wire  io_c2b_rst_reg_io_q; // @[AsyncResetReg.scala 74:21]
  wire  io_c2b_rst_reg_io_clk; // @[AsyncResetReg.scala 74:21]
  wire  io_c2b_rst_reg_io_rst; // @[AsyncResetReg.scala 74:21]
  reg [19:0] rx_a; // @[TX.scala 31:19]
  reg [19:0] rx_b; // @[TX.scala 31:19]
  reg [19:0] rx_c; // @[TX.scala 31:19]
  reg [19:0] rx_d; // @[TX.scala 31:19]
  reg [19:0] rx_e; // @[TX.scala 31:19]
  reg [19:0] tx_a; // @[TX.scala 32:19]
  reg [19:0] tx_b; // @[TX.scala 32:19]
  reg [19:0] tx_c; // @[TX.scala 32:19]
  reg [19:0] tx_d; // @[TX.scala 32:19]
  reg [19:0] tx_e; // @[TX.scala 32:19]
  wire  _ioX_first_T = qa_q_io_deq_ready & qa_q_io_deq_valid; // @[Decoupled.scala 40:37]
  reg  ioX_first; // @[Reg.scala 27:20]
  wire  _GEN_0 = _ioX_first_T ? qa_q_io_deq_bits_last : ioX_first; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [19:0] _GEN_19 = {{13'd0}, qa_q_io_deq_bits_beats}; // @[TX.scala 52:24]
  wire [20:0] ioX_delta = tx_a - _GEN_19; // @[TX.scala 52:24]
  wire [20:0] _ioX_allow_T_1 = tx_a - _GEN_19; // @[TX.scala 53:34]
  wire  ioX_allow = ~ioX_first | $signed(_ioX_allow_T_1) >= 21'sh0; // @[TX.scala 53:24]
  wire [20:0] _ioX_tx_a_T_2 = _ioX_first_T & ioX_first ? ioX_delta : {{1'd0}, tx_a}; // @[TX.scala 54:18]
  wire  _ioX_tx_a_T_3 = txInc_sink_io_deq_ready & txInc_sink_io_deq_valid; // @[Decoupled.scala 40:37]
  wire [19:0] _ioX_tx_a_T_4 = _ioX_tx_a_T_3 ? txInc_sink_io_deq_bits_a : 20'h0; // @[TX.scala 54:58]
  wire [20:0] _GEN_20 = {{1'd0}, _ioX_tx_a_T_4}; // @[TX.scala 54:53]
  wire [20:0] _ioX_tx_a_T_6 = _ioX_tx_a_T_2 + _GEN_20; // @[TX.scala 54:53]
  wire  _ioX_first_T_1 = qb_q_io_deq_ready & qb_q_io_deq_valid; // @[Decoupled.scala 40:37]
  reg  ioX_first_1; // @[Reg.scala 27:20]
  wire  _GEN_1 = _ioX_first_T_1 ? qb_q_io_deq_bits_last : ioX_first_1; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [19:0] _GEN_21 = {{13'd0}, qb_q_io_deq_bits_beats}; // @[TX.scala 52:24]
  wire [20:0] ioX_delta_1 = tx_b - _GEN_21; // @[TX.scala 52:24]
  wire [20:0] _ioX_allow_T_4 = tx_b - _GEN_21; // @[TX.scala 53:34]
  wire  ioX_allow_1 = ~ioX_first_1 | $signed(_ioX_allow_T_4) >= 21'sh0; // @[TX.scala 53:24]
  wire [20:0] _ioX_tx_bT_2 = _ioX_first_T_1 & ioX_first_1 ? ioX_delta_1 : {{1'd0}, tx_b}; // @[TX.scala 54:18]
  wire [19:0] _ioX_tx_bT_4 = _ioX_tx_a_T_3 ? txInc_sink_io_deq_bits_b : 20'h0; // @[TX.scala 54:58]
  wire [20:0] _GEN_22 = {{1'd0}, _ioX_tx_bT_4}; // @[TX.scala 54:53]
  wire [20:0] _ioX_tx_bT_6 = _ioX_tx_bT_2 + _GEN_22; // @[TX.scala 54:53]
  wire  _ioX_first_T_2 = qc_q_io_deq_ready & qc_q_io_deq_valid; // @[Decoupled.scala 40:37]
  reg  ioX_first_2; // @[Reg.scala 27:20]
  wire  _GEN_2 = _ioX_first_T_2 ? qc_q_io_deq_bits_last : ioX_first_2; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [19:0] _GEN_23 = {{13'd0}, qc_q_io_deq_bits_beats}; // @[TX.scala 52:24]
  wire [20:0] ioX_delta_2 = tx_c - _GEN_23; // @[TX.scala 52:24]
  wire [20:0] _ioX_allow_T_7 = tx_c - _GEN_23; // @[TX.scala 53:34]
  wire  ioX_allow_2 = ~ioX_first_2 | $signed(_ioX_allow_T_7) >= 21'sh0; // @[TX.scala 53:24]
  wire [20:0] _ioX_tx_c_T_2 = _ioX_first_T_2 & ioX_first_2 ? ioX_delta_2 : {{1'd0}, tx_c}; // @[TX.scala 54:18]
  wire [19:0] _ioX_tx_c_T_4 = _ioX_tx_a_T_3 ? txInc_sink_io_deq_bits_c : 20'h0; // @[TX.scala 54:58]
  wire [20:0] _GEN_24 = {{1'd0}, _ioX_tx_c_T_4}; // @[TX.scala 54:53]
  wire [20:0] _ioX_tx_c_T_6 = _ioX_tx_c_T_2 + _GEN_24; // @[TX.scala 54:53]
  wire  _ioX_first_T_3 = qd_q_io_deq_ready & qd_q_io_deq_valid; // @[Decoupled.scala 40:37]
  reg  ioX_first_3; // @[Reg.scala 27:20]
  wire  _GEN_3 = _ioX_first_T_3 ? qd_q_io_deq_bits_last : ioX_first_3; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [19:0] _GEN_25 = {{13'd0}, qd_q_io_deq_bits_beats}; // @[TX.scala 52:24]
  wire [20:0] ioX_delta_3 = tx_d - _GEN_25; // @[TX.scala 52:24]
  wire [20:0] _ioX_allow_T_10 = tx_d - _GEN_25; // @[TX.scala 53:34]
  wire  ioX_allow_3 = ~ioX_first_3 | $signed(_ioX_allow_T_10) >= 21'sh0; // @[TX.scala 53:24]
  wire [20:0] _ioX_tx_d_T_2 = _ioX_first_T_3 & ioX_first_3 ? ioX_delta_3 : {{1'd0}, tx_d}; // @[TX.scala 54:18]
  wire [19:0] _ioX_tx_d_T_4 = _ioX_tx_a_T_3 ? txInc_sink_io_deq_bits_d : 20'h0; // @[TX.scala 54:58]
  wire [20:0] _GEN_26 = {{1'd0}, _ioX_tx_d_T_4}; // @[TX.scala 54:53]
  wire [20:0] _ioX_tx_d_T_6 = _ioX_tx_d_T_2 + _GEN_26; // @[TX.scala 54:53]
  wire  _ioX_first_T_4 = qe_q_io_deq_ready & qe_q_io_deq_valid; // @[Decoupled.scala 40:37]
  reg  ioX_first_4; // @[Reg.scala 27:20]
  wire  _GEN_4 = _ioX_first_T_4 ? qe_q_io_deq_bits_last : ioX_first_4; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [19:0] _GEN_27 = {{13'd0}, qe_q_io_deq_bits_beats}; // @[TX.scala 52:24]
  wire [20:0] ioX_delta_4 = tx_e - _GEN_27; // @[TX.scala 52:24]
  wire [20:0] _ioX_allow_T_13 = tx_e - _GEN_27; // @[TX.scala 53:34]
  wire  ioX_allow_4 = ~ioX_first_4 | $signed(_ioX_allow_T_13) >= 21'sh0; // @[TX.scala 53:24]
  wire [20:0] _ioX_tx_e_T_2 = _ioX_first_T_4 & ioX_first_4 ? ioX_delta_4 : {{1'd0}, tx_e}; // @[TX.scala 54:18]
  wire [19:0] _ioX_tx_e_T_4 = _ioX_tx_a_T_3 ? txInc_sink_io_deq_bits_e : 20'h0; // @[TX.scala 54:58]
  wire [20:0] _GEN_28 = {{1'd0}, _ioX_tx_e_T_4}; // @[TX.scala 54:53]
  wire [20:0] _ioX_tx_e_T_6 = _ioX_tx_e_T_2 + _GEN_28; // @[TX.scala 54:53]
  wire [19:0] _GEN_29 = {{1'd0}, rx_a[19:1]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_1 = rx_a | _GEN_29; // @[package.scala 253:43]
  wire [19:0] _GEN_30 = {{2'd0}, _mask_T_1[19:2]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_3 = _mask_T_1 | _GEN_30; // @[package.scala 253:43]
  wire [19:0] _GEN_31 = {{4'd0}, _mask_T_3[19:4]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_5 = _mask_T_3 | _GEN_31; // @[package.scala 253:43]
  wire [19:0] _GEN_32 = {{8'd0}, _mask_T_5[19:8]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_7 = _mask_T_5 | _GEN_32; // @[package.scala 253:43]
  wire [19:0] _GEN_33 = {{16'd0}, _mask_T_7[19:16]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_9 = _mask_T_7 | _GEN_33; // @[package.scala 253:43]
  wire [18:0] mask = _mask_T_9[19:1]; // @[Bundles.scala 47:29]
  wire [19:0] _msbOH_T = ~rx_a; // @[Bundles.scala 48:21]
  wire [19:0] _GEN_34 = {{1'd0}, mask}; // @[Bundles.scala 48:24]
  wire [19:0] _msbOH_T_1 = _msbOH_T | _GEN_34; // @[Bundles.scala 48:24]
  wire [19:0] msbOH = ~_msbOH_T_1; // @[Bundles.scala 48:19]
  wire [20:0] _msb_T = {msbOH, 1'h0}; // @[Bundles.scala 49:32]
  wire [4:0] msb_hi = _msb_T[20:16]; // @[OneHot.scala 30:18]
  wire [15:0] msb_lo = _msb_T[15:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_1 = |msb_hi; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_35 = {{11'd0}, msb_hi}; // @[OneHot.scala 32:28]
  wire [15:0] _msb_T_1 = _GEN_35 | msb_lo; // @[OneHot.scala 32:28]
  wire [7:0] msb_hi_2 = _msb_T_1[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] msb_lo_1 = _msb_T_1[7:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_3 = |msb_hi_2; // @[OneHot.scala 32:14]
  wire [7:0] _msb_T_2 = msb_hi_2 | msb_lo_1; // @[OneHot.scala 32:28]
  wire [3:0] msb_hi_4 = _msb_T_2[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] msb_lo_2 = _msb_T_2[3:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_5 = |msb_hi_4; // @[OneHot.scala 32:14]
  wire [3:0] _msb_T_3 = msb_hi_4 | msb_lo_2; // @[OneHot.scala 32:28]
  wire [1:0] msb_hi_6 = _msb_T_3[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] msb_lo_3 = _msb_T_3[1:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_7 = |msb_hi_6; // @[OneHot.scala 32:14]
  wire [1:0] _msb_T_4 = msb_hi_6 | msb_lo_3; // @[OneHot.scala 32:28]
  wire  msb_lo_4 = _msb_T_4[1]; // @[CircuitMath.scala 30:8]
  wire [19:0] a_rest = rx_a & _GEN_34; // @[Bundles.scala 51:15]
  wire [19:0] _GEN_37 = {{1'd0}, rx_b[19:1]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_12 = rx_b | _GEN_37; // @[package.scala 253:43]
  wire [19:0] _GEN_38 = {{2'd0}, _mask_T_12[19:2]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_14 = _mask_T_12 | _GEN_38; // @[package.scala 253:43]
  wire [19:0] _GEN_39 = {{4'd0}, _mask_T_14[19:4]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_16 = _mask_T_14 | _GEN_39; // @[package.scala 253:43]
  wire [19:0] _GEN_40 = {{8'd0}, _mask_T_16[19:8]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_18 = _mask_T_16 | _GEN_40; // @[package.scala 253:43]
  wire [19:0] _GEN_41 = {{16'd0}, _mask_T_18[19:16]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_20 = _mask_T_18 | _GEN_41; // @[package.scala 253:43]
  wire [18:0] mask_1 = _mask_T_20[19:1]; // @[Bundles.scala 47:29]
  wire [19:0] _msbOH_T_2 = ~rx_b; // @[Bundles.scala 48:21]
  wire [19:0] _GEN_42 = {{1'd0}, mask_1}; // @[Bundles.scala 48:24]
  wire [19:0] _msbOH_T_3 = _msbOH_T_2 | _GEN_42; // @[Bundles.scala 48:24]
  wire [19:0] msbOH_1 = ~_msbOH_T_3; // @[Bundles.scala 48:19]
  wire [20:0] _msb_T_5 = {msbOH_1, 1'h0}; // @[Bundles.scala 49:32]
  wire [4:0] msb_hi_8 = _msb_T_5[20:16]; // @[OneHot.scala 30:18]
  wire [15:0] msb_lo_8 = _msb_T_5[15:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_9 = |msb_hi_8; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_43 = {{11'd0}, msb_hi_8}; // @[OneHot.scala 32:28]
  wire [15:0] _msb_T_6 = _GEN_43 | msb_lo_8; // @[OneHot.scala 32:28]
  wire [7:0] msb_hi_10 = _msb_T_6[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] msb_lo_9 = _msb_T_6[7:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_11 = |msb_hi_10; // @[OneHot.scala 32:14]
  wire [7:0] _msb_T_7 = msb_hi_10 | msb_lo_9; // @[OneHot.scala 32:28]
  wire [3:0] msb_hi_12 = _msb_T_7[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] msb_lo_10 = _msb_T_7[3:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_13 = |msb_hi_12; // @[OneHot.scala 32:14]
  wire [3:0] _msb_T_8 = msb_hi_12 | msb_lo_10; // @[OneHot.scala 32:28]
  wire [1:0] msb_hi_14 = _msb_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] msb_lo_11 = _msb_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_15 = |msb_hi_14; // @[OneHot.scala 32:14]
  wire [1:0] _msb_T_9 = msb_hi_14 | msb_lo_11; // @[OneHot.scala 32:28]
  wire  msb_lo_12 = _msb_T_9[1]; // @[CircuitMath.scala 30:8]
  wire [19:0] b_rest = rx_b & _GEN_42; // @[Bundles.scala 51:15]
  wire [19:0] _GEN_45 = {{1'd0}, rx_c[19:1]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_23 = rx_c | _GEN_45; // @[package.scala 253:43]
  wire [19:0] _GEN_46 = {{2'd0}, _mask_T_23[19:2]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_25 = _mask_T_23 | _GEN_46; // @[package.scala 253:43]
  wire [19:0] _GEN_47 = {{4'd0}, _mask_T_25[19:4]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_27 = _mask_T_25 | _GEN_47; // @[package.scala 253:43]
  wire [19:0] _GEN_48 = {{8'd0}, _mask_T_27[19:8]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_29 = _mask_T_27 | _GEN_48; // @[package.scala 253:43]
  wire [19:0] _GEN_49 = {{16'd0}, _mask_T_29[19:16]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_31 = _mask_T_29 | _GEN_49; // @[package.scala 253:43]
  wire [18:0] mask_2 = _mask_T_31[19:1]; // @[Bundles.scala 47:29]
  wire [19:0] _msbOH_T_4 = ~rx_c; // @[Bundles.scala 48:21]
  wire [19:0] _GEN_50 = {{1'd0}, mask_2}; // @[Bundles.scala 48:24]
  wire [19:0] _msbOH_T_5 = _msbOH_T_4 | _GEN_50; // @[Bundles.scala 48:24]
  wire [19:0] msbOH_2 = ~_msbOH_T_5; // @[Bundles.scala 48:19]
  wire [20:0] _msb_T_10 = {msbOH_2, 1'h0}; // @[Bundles.scala 49:32]
  wire [4:0] msb_hi_16 = _msb_T_10[20:16]; // @[OneHot.scala 30:18]
  wire [15:0] msb_lo_16 = _msb_T_10[15:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_17 = |msb_hi_16; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_51 = {{11'd0}, msb_hi_16}; // @[OneHot.scala 32:28]
  wire [15:0] _msb_T_11 = _GEN_51 | msb_lo_16; // @[OneHot.scala 32:28]
  wire [7:0] msb_hi_18 = _msb_T_11[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] msb_lo_17 = _msb_T_11[7:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_19 = |msb_hi_18; // @[OneHot.scala 32:14]
  wire [7:0] _msb_T_12 = msb_hi_18 | msb_lo_17; // @[OneHot.scala 32:28]
  wire [3:0] msb_hi_20 = _msb_T_12[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] msb_lo_18 = _msb_T_12[3:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_21 = |msb_hi_20; // @[OneHot.scala 32:14]
  wire [3:0] _msb_T_13 = msb_hi_20 | msb_lo_18; // @[OneHot.scala 32:28]
  wire [1:0] msb_hi_22 = _msb_T_13[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] msb_lo_19 = _msb_T_13[1:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_23 = |msb_hi_22; // @[OneHot.scala 32:14]
  wire [1:0] _msb_T_14 = msb_hi_22 | msb_lo_19; // @[OneHot.scala 32:28]
  wire  msb_lo_20 = _msb_T_14[1]; // @[CircuitMath.scala 30:8]
  wire [19:0] c_rest = rx_c & _GEN_50; // @[Bundles.scala 51:15]
  wire [19:0] _GEN_53 = {{1'd0}, rx_d[19:1]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_34 = rx_d | _GEN_53; // @[package.scala 253:43]
  wire [19:0] _GEN_54 = {{2'd0}, _mask_T_34[19:2]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_36 = _mask_T_34 | _GEN_54; // @[package.scala 253:43]
  wire [19:0] _GEN_55 = {{4'd0}, _mask_T_36[19:4]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_38 = _mask_T_36 | _GEN_55; // @[package.scala 253:43]
  wire [19:0] _GEN_56 = {{8'd0}, _mask_T_38[19:8]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_40 = _mask_T_38 | _GEN_56; // @[package.scala 253:43]
  wire [19:0] _GEN_57 = {{16'd0}, _mask_T_40[19:16]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_42 = _mask_T_40 | _GEN_57; // @[package.scala 253:43]
  wire [18:0] mask_3 = _mask_T_42[19:1]; // @[Bundles.scala 47:29]
  wire [19:0] _msbOH_T_6 = ~rx_d; // @[Bundles.scala 48:21]
  wire [19:0] _GEN_58 = {{1'd0}, mask_3}; // @[Bundles.scala 48:24]
  wire [19:0] _msbOH_T_7 = _msbOH_T_6 | _GEN_58; // @[Bundles.scala 48:24]
  wire [19:0] msbOH_3 = ~_msbOH_T_7; // @[Bundles.scala 48:19]
  wire [20:0] _msb_T_15 = {msbOH_3, 1'h0}; // @[Bundles.scala 49:32]
  wire [4:0] msb_hi_24 = _msb_T_15[20:16]; // @[OneHot.scala 30:18]
  wire [15:0] msb_lo_24 = _msb_T_15[15:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_25 = |msb_hi_24; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_59 = {{11'd0}, msb_hi_24}; // @[OneHot.scala 32:28]
  wire [15:0] _msb_T_16 = _GEN_59 | msb_lo_24; // @[OneHot.scala 32:28]
  wire [7:0] msb_hi_26 = _msb_T_16[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] msb_lo_25 = _msb_T_16[7:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_27 = |msb_hi_26; // @[OneHot.scala 32:14]
  wire [7:0] _msb_T_17 = msb_hi_26 | msb_lo_25; // @[OneHot.scala 32:28]
  wire [3:0] msb_hi_28 = _msb_T_17[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] msb_lo_26 = _msb_T_17[3:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_29 = |msb_hi_28; // @[OneHot.scala 32:14]
  wire [3:0] _msb_T_18 = msb_hi_28 | msb_lo_26; // @[OneHot.scala 32:28]
  wire [1:0] msb_hi_30 = _msb_T_18[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] msb_lo_27 = _msb_T_18[1:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_31 = |msb_hi_30; // @[OneHot.scala 32:14]
  wire [1:0] _msb_T_19 = msb_hi_30 | msb_lo_27; // @[OneHot.scala 32:28]
  wire  msb_lo_28 = _msb_T_19[1]; // @[CircuitMath.scala 30:8]
  wire [19:0] d_rest = rx_d & _GEN_58; // @[Bundles.scala 51:15]
  wire [19:0] _GEN_61 = {{1'd0}, rx_e[19:1]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_45 = rx_e | _GEN_61; // @[package.scala 253:43]
  wire [19:0] _GEN_62 = {{2'd0}, _mask_T_45[19:2]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_47 = _mask_T_45 | _GEN_62; // @[package.scala 253:43]
  wire [19:0] _GEN_63 = {{4'd0}, _mask_T_47[19:4]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_49 = _mask_T_47 | _GEN_63; // @[package.scala 253:43]
  wire [19:0] _GEN_64 = {{8'd0}, _mask_T_49[19:8]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_51 = _mask_T_49 | _GEN_64; // @[package.scala 253:43]
  wire [19:0] _GEN_65 = {{16'd0}, _mask_T_51[19:16]}; // @[package.scala 253:43]
  wire [19:0] _mask_T_53 = _mask_T_51 | _GEN_65; // @[package.scala 253:43]
  wire [18:0] mask_4 = _mask_T_53[19:1]; // @[Bundles.scala 47:29]
  wire [19:0] _msbOH_T_8 = ~rx_e; // @[Bundles.scala 48:21]
  wire [19:0] _GEN_66 = {{1'd0}, mask_4}; // @[Bundles.scala 48:24]
  wire [19:0] _msbOH_T_9 = _msbOH_T_8 | _GEN_66; // @[Bundles.scala 48:24]
  wire [19:0] msbOH_4 = ~_msbOH_T_9; // @[Bundles.scala 48:19]
  wire [20:0] _msb_T_20 = {msbOH_4, 1'h0}; // @[Bundles.scala 49:32]
  wire [4:0] msb_hi_32 = _msb_T_20[20:16]; // @[OneHot.scala 30:18]
  wire [15:0] msb_lo_32 = _msb_T_20[15:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_33 = |msb_hi_32; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_67 = {{11'd0}, msb_hi_32}; // @[OneHot.scala 32:28]
  wire [15:0] _msb_T_21 = _GEN_67 | msb_lo_32; // @[OneHot.scala 32:28]
  wire [7:0] msb_hi_34 = _msb_T_21[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] msb_lo_33 = _msb_T_21[7:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_35 = |msb_hi_34; // @[OneHot.scala 32:14]
  wire [7:0] _msb_T_22 = msb_hi_34 | msb_lo_33; // @[OneHot.scala 32:28]
  wire [3:0] msb_hi_36 = _msb_T_22[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] msb_lo_34 = _msb_T_22[3:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_37 = |msb_hi_36; // @[OneHot.scala 32:14]
  wire [3:0] _msb_T_23 = msb_hi_36 | msb_lo_34; // @[OneHot.scala 32:28]
  wire [1:0] msb_hi_38 = _msb_T_23[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] msb_lo_35 = _msb_T_23[1:0]; // @[OneHot.scala 31:18]
  wire  msb_hi_39 = |msb_hi_38; // @[OneHot.scala 32:14]
  wire [1:0] _msb_T_24 = msb_hi_38 | msb_lo_35; // @[OneHot.scala 32:28]
  wire  msb_lo_36 = _msb_T_24[1]; // @[CircuitMath.scala 30:8]
  wire [19:0] e_rest = rx_e & _GEN_66; // @[Bundles.scala 51:15]
  wire [11:0] header_lo = {msb_hi_1,msb_hi_3,msb_hi_5,msb_hi_7,msb_lo_4,4'h0,3'h5}; // @[Cat.scala 30:58]
  wire [9:0] header_hi_lo = {msb_hi_17,msb_hi_19,msb_hi_21,msb_hi_23,msb_lo_20,msb_hi_9,msb_hi_11,msb_hi_13,msb_hi_15,
    msb_lo_12}; // @[Cat.scala 30:58]
  wire [9:0] header_hi_hi = {msb_hi_33,msb_hi_35,msb_hi_37,msb_hi_39,msb_lo_36,msb_hi_25,msb_hi_27,msb_hi_29,msb_hi_31,
    msb_lo_28}; // @[Cat.scala 30:58]
  wire [19:0] header_hi = {header_hi_hi,header_hi_lo}; // @[Cat.scala 30:58]
  wire [31:0] rxHeader = {header_hi_hi,header_hi_lo,msb_hi_1,msb_hi_3,msb_hi_5,msb_hi_7,msb_lo_4,4'h0,3'h5}; // @[Cat.scala 30:58]
  wire  _rx_T = rxQ_io_enq_ready & rxQ_io_enq_valid; // @[Decoupled.scala 40:37]
  wire [19:0] _rx_T_1_a = _rx_T ? a_rest : rx_a; // @[TX.scala 70:12]
  wire [19:0] _rx_T_1_b = _rx_T ? b_rest : rx_b; // @[TX.scala 70:12]
  wire [19:0] _rx_T_1_c = _rx_T ? c_rest : rx_c; // @[TX.scala 70:12]
  wire [19:0] _rx_T_1_d = _rx_T ? d_rest : rx_d; // @[TX.scala 70:12]
  wire [19:0] _rx_T_1_e = _rx_T ? e_rest : rx_e; // @[TX.scala 70:12]
  wire  _rx_T_2 = rxInc_sink_io_deq_ready & rxInc_sink_io_deq_valid; // @[Decoupled.scala 40:37]
  wire [19:0] _rx_T_3_a = _rx_T_2 ? rxInc_sink_io_deq_bits_a : 20'h0; // @[TX.scala 70:49]
  wire [19:0] _rx_T_3_b = _rx_T_2 ? rxInc_sink_io_deq_bits_b : 20'h0; // @[TX.scala 70:49]
  wire [19:0] _rx_T_3_c = _rx_T_2 ? rxInc_sink_io_deq_bits_c : 20'h0; // @[TX.scala 70:49]
  wire [19:0] _rx_T_3_d = _rx_T_2 ? rxInc_sink_io_deq_bits_d : 20'h0; // @[TX.scala 70:49]
  wire [19:0] _rx_T_3_e = _rx_T_2 ? rxInc_sink_io_deq_bits_e : 20'h0; // @[TX.scala 70:49]
  wire [20:0] rx_z = _rx_T_1_a + _rx_T_3_a; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_a_T_3 = |rx_z[20] ? 21'hfffff : rx_z; // @[Bundles.scala 39:15]
  wire [20:0] rx_z_1 = _rx_T_1_b + _rx_T_3_b; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_bT_3 = |rx_z_1[20] ? 21'hfffff : rx_z_1; // @[Bundles.scala 39:15]
  wire [20:0] rx_z_2 = _rx_T_1_c + _rx_T_3_c; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_c_T_3 = |rx_z_2[20] ? 21'hfffff : rx_z_2; // @[Bundles.scala 39:15]
  wire [20:0] rx_z_3 = _rx_T_1_d + _rx_T_3_d; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_d_T_3 = |rx_z_3[20] ? 21'hfffff : rx_z_3; // @[Bundles.scala 39:15]
  wire [20:0] rx_z_4 = _rx_T_1_e + _rx_T_3_e; // @[Bundles.scala 38:17]
  wire [20:0] _rx_out_e_T_3 = |rx_z_4[20] ? 21'hfffff : rx_z_4; // @[Bundles.scala 39:15]
  reg [1:0] xmit; // @[TX.scala 80:21]
  wire  forceXmit = xmit == 2'h0; // @[TX.scala 81:24]
  wire  allowReturn = ~(ioX_cq_io_deq_valid | ioX_cq_1_io_deq_valid | ioX_cq_2_io_deq_valid | ioX_cq_3_io_deq_valid |
    ioX_cq_4_io_deq_valid) | forceXmit; // @[TX.scala 86:54]
  wire  f_valid = rxQ_io_deq_valid & allowReturn; // @[TX.scala 88:31]
  wire [5:0] requests = {f_valid,ioX_cq_4_io_deq_valid,ioX_cq_3_io_deq_valid,ioX_cq_2_io_deq_valid,ioX_cq_1_io_deq_valid
    ,ioX_cq_io_deq_valid}; // @[Cat.scala 30:58]
  wire  f_bits_last = rxQ_io_deq_bits_last; // @[TX.scala 73:15 TX.scala 87:11]
  wire [5:0] lasts = {f_bits_last,ioX_cq_4_io_deq_bits_last,ioX_cq_3_io_deq_bits_last,ioX_cq_2_io_deq_bits_last,
    ioX_cq_1_io_deq_bits_last,ioX_cq_io_deq_bits_last}; // @[Cat.scala 30:58]
  wire [1:0] _xmit_T_1 = xmit - 2'h1; // @[TX.scala 82:36]
  reg  first; // @[TX.scala 92:22]
  reg [5:0] readys_mask; // @[Arbiter.scala 23:23]
  wire [5:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 24:30]
  wire [5:0] readys_filter_hi = requests & _readys_filter_T; // @[Arbiter.scala 24:28]
  wire [11:0] readys_filter = {readys_filter_hi,f_valid,ioX_cq_4_io_deq_valid,ioX_cq_3_io_deq_valid,
    ioX_cq_2_io_deq_valid,ioX_cq_1_io_deq_valid,ioX_cq_io_deq_valid}; // @[Cat.scala 30:58]
  wire [11:0] _GEN_69 = {{1'd0}, readys_filter[11:1]}; // @[package.scala 253:43]
  wire [11:0] _readys_unready_T_1 = readys_filter | _GEN_69; // @[package.scala 253:43]
  wire [11:0] _GEN_70 = {{2'd0}, _readys_unready_T_1[11:2]}; // @[package.scala 253:43]
  wire [11:0] _readys_unready_T_3 = _readys_unready_T_1 | _GEN_70; // @[package.scala 253:43]
  wire [11:0] _GEN_71 = {{4'd0}, _readys_unready_T_3[11:4]}; // @[package.scala 253:43]
  wire [11:0] _readys_unready_T_5 = _readys_unready_T_3 | _GEN_71; // @[package.scala 253:43]
  wire [11:0] _readys_unready_T_8 = {readys_mask, 6'h0}; // @[Arbiter.scala 25:66]
  wire [11:0] _GEN_72 = {{1'd0}, _readys_unready_T_5[11:1]}; // @[Arbiter.scala 25:58]
  wire [11:0] readys_unready = _GEN_72 | _readys_unready_T_8; // @[Arbiter.scala 25:58]
  wire [5:0] _readys_readys_T_2 = readys_unready[11:6] & readys_unready[5:0]; // @[Arbiter.scala 26:39]
  wire [5:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  reg [5:0] state; // @[TX.scala 93:18]
  wire [5:0] allowed = first ? readys_readys : state; // @[TX.scala 97:20]
  reg  txBusy; // @[TX.scala 99:23]
  wire  f_ready = allowed[5] & ~txBusy; // @[TX.scala 100:77]
  wire  _T_1 = f_ready & f_valid; // @[Decoupled.scala 40:37]
  wire [5:0] _readys_mask_T = readys_readys & requests; // @[Arbiter.scala 28:29]
  wire [6:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  wire [5:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[5:0]; // @[package.scala 244:43]
  wire [7:0] _readys_mask_T_4 = {_readys_mask_T_3, 2'h0}; // @[package.scala 244:48]
  wire [5:0] _readys_mask_T_6 = _readys_mask_T_3 | _readys_mask_T_4[5:0]; // @[package.scala 244:43]
  wire [9:0] _readys_mask_T_7 = {_readys_mask_T_6, 4'h0}; // @[package.scala 244:48]
  wire [5:0] _readys_mask_T_9 = _readys_mask_T_6 | _readys_mask_T_7[5:0]; // @[package.scala 244:43]
  wire [5:0] grant = first ? _readys_mask_T : state; // @[TX.scala 96:18]
  wire  _send_T = ioX_cq_io_deq_ready & ioX_cq_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _send_T_1 = ioX_cq_1_io_deq_ready & ioX_cq_1_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _send_T_2 = ioX_cq_2_io_deq_ready & ioX_cq_2_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _send_T_3 = ioX_cq_3_io_deq_ready & ioX_cq_3_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _send_T_4 = ioX_cq_4_io_deq_ready & ioX_cq_4_io_deq_valid; // @[Decoupled.scala 40:37]
  wire  send = _send_T | _send_T_1 | _send_T_2 | _send_T_3 | _send_T_4 | _T_1; // @[package.scala 72:59]
  wire [5:0] _first_T = grant & lasts; // @[TX.scala 105:33]
  wire  _GEN_8 = send ? |_first_T : first; // @[TX.scala 105:15 TX.scala 105:23 TX.scala 92:22]
  reg [1:0] transferByteCnt; // @[TX.scala 108:32]
  wire  _GEN_10 = send | txBusy; // @[TX.scala 109:14 TX.scala 110:12 TX.scala 99:23]
  wire [1:0] _transferByteCnt_T_1 = transferByteCnt + 2'h1; // @[TX.scala 113:40]
  wire [31:0] _transferDataReg_WIRE__0 = ioX_cq_io_deq_bits_data; // @[TX.scala 118:51 TX.scala 118:51]
  wire [31:0] _transferDataReg_T_6 = grant[0] ? _transferDataReg_WIRE__0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_WIRE__1 = ioX_cq_1_io_deq_bits_data; // @[TX.scala 118:51 TX.scala 118:51]
  wire [31:0] _transferDataReg_T_7 = grant[1] ? _transferDataReg_WIRE__1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_WIRE__2 = ioX_cq_2_io_deq_bits_data; // @[TX.scala 118:51 TX.scala 118:51]
  wire [31:0] _transferDataReg_T_8 = grant[2] ? _transferDataReg_WIRE__2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_WIRE__3 = ioX_cq_3_io_deq_bits_data; // @[TX.scala 118:51 TX.scala 118:51]
  wire [31:0] _transferDataReg_T_9 = grant[3] ? _transferDataReg_WIRE__3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_WIRE__4 = ioX_cq_4_io_deq_bits_data; // @[TX.scala 118:51 TX.scala 118:51]
  wire [31:0] _transferDataReg_T_10 = grant[4] ? _transferDataReg_WIRE__4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] f_bits_data = rxQ_io_deq_bits_data; // @[TX.scala 73:15 TX.scala 87:11]
  wire [31:0] _transferDataReg_T_11 = grant[5] ? f_bits_data : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_T_12 = _transferDataReg_T_6 | _transferDataReg_T_7; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_T_13 = _transferDataReg_T_12 | _transferDataReg_T_8; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_T_14 = _transferDataReg_T_13 | _transferDataReg_T_9; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_T_15 = _transferDataReg_T_14 | _transferDataReg_T_10; // @[Mux.scala 27:72]
  wire [31:0] _transferDataReg_T_16 = _transferDataReg_T_15 | _transferDataReg_T_11; // @[Mux.scala 27:72]
  reg [31:0] transferDataReg; // @[Reg.scala 15:16]
  wire [7:0] transferBytes_0 = transferDataReg[31:24]; // @[TX.scala 119:42]
  wire [7:0] transferBytes_1 = transferDataReg[23:16]; // @[TX.scala 119:67]
  wire [7:0] transferBytes_2 = transferDataReg[15:8]; // @[TX.scala 119:92]
  wire [7:0] transferBytes_3 = transferDataReg[7:0]; // @[TX.scala 119:116]
  reg  io_c2b_send_REG; // @[TX.scala 124:33]
  reg  io_c2b_send_REG_1; // @[TX.scala 124:25]
  reg [7:0] io_c2b_data_REG; // @[TX.scala 125:33]
  reg [7:0] io_c2b_data_REG_1; // @[TX.scala 125:25]
  wire [19:0] rx_out_2_a = _rx_out_a_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] rx_out_2_b = _rx_out_bT_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] rx_out_2_c = _rx_out_c_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] rx_out_2_d = _rx_out_d_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  wire [19:0] rx_out_2_e = _rx_out_e_T_3[19:0]; // @[Bundles.scala 36:19 Bundles.scala 39:9]
  AsyncQueueSink_5 rxInc_sink ( // @[AsyncQueue.scala 207:22]
    .clock(rxInc_sink_clock),
    .reset(rxInc_sink_reset),
    .io_deq_ready(rxInc_sink_io_deq_ready),
    .io_deq_valid(rxInc_sink_io_deq_valid),
    .io_deq_bits_a(rxInc_sink_io_deq_bits_a),
    .io_deq_bits_b(rxInc_sink_io_deq_bits_b),
    .io_deq_bits_c(rxInc_sink_io_deq_bits_c),
    .io_deq_bits_d(rxInc_sink_io_deq_bits_d),
    .io_deq_bits_e(rxInc_sink_io_deq_bits_e),
    .io_async_mem_0_a(rxInc_sink_io_async_mem_0_a),
    .io_async_mem_0_b(rxInc_sink_io_async_mem_0_b),
    .io_async_mem_0_c(rxInc_sink_io_async_mem_0_c),
    .io_async_mem_0_d(rxInc_sink_io_async_mem_0_d),
    .io_async_mem_0_e(rxInc_sink_io_async_mem_0_e),
    .io_async_ridx(rxInc_sink_io_async_ridx),
    .io_async_widx(rxInc_sink_io_async_widx),
    .io_async_safe_ridx_valid(rxInc_sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(rxInc_sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(rxInc_sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(rxInc_sink_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink_5 txInc_sink ( // @[AsyncQueue.scala 207:22]
    .clock(txInc_sink_clock),
    .reset(txInc_sink_reset),
    .io_deq_ready(txInc_sink_io_deq_ready),
    .io_deq_valid(txInc_sink_io_deq_valid),
    .io_deq_bits_a(txInc_sink_io_deq_bits_a),
    .io_deq_bits_b(txInc_sink_io_deq_bits_b),
    .io_deq_bits_c(txInc_sink_io_deq_bits_c),
    .io_deq_bits_d(txInc_sink_io_deq_bits_d),
    .io_deq_bits_e(txInc_sink_io_deq_bits_e),
    .io_async_mem_0_a(txInc_sink_io_async_mem_0_a),
    .io_async_mem_0_b(txInc_sink_io_async_mem_0_b),
    .io_async_mem_0_c(txInc_sink_io_async_mem_0_c),
    .io_async_mem_0_d(txInc_sink_io_async_mem_0_d),
    .io_async_mem_0_e(txInc_sink_io_async_mem_0_e),
    .io_async_ridx(txInc_sink_io_async_ridx),
    .io_async_widx(txInc_sink_io_async_widx),
    .io_async_safe_ridx_valid(txInc_sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(txInc_sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(txInc_sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(txInc_sink_io_async_safe_sink_reset_n)
  );
  ShiftQueue qa_q ( // @[ShiftQueue.scala 60:19]
    .clock(qa_q_clock),
    .reset(qa_q_reset),
    .io_enq_ready(qa_q_io_enq_ready),
    .io_enq_valid(qa_q_io_enq_valid),
    .io_enq_bits_data(qa_q_io_enq_bits_data),
    .io_enq_bits_last(qa_q_io_enq_bits_last),
    .io_enq_bits_beats(qa_q_io_enq_bits_beats),
    .io_deq_ready(qa_q_io_deq_ready),
    .io_deq_valid(qa_q_io_deq_valid),
    .io_deq_bits_data(qa_q_io_deq_bits_data),
    .io_deq_bits_last(qa_q_io_deq_bits_last),
    .io_deq_bits_beats(qa_q_io_deq_bits_beats)
  );
  ShiftQueue qb_q ( // @[ShiftQueue.scala 60:19]
    .clock(qb_q_clock),
    .reset(qb_q_reset),
    .io_enq_ready(qb_q_io_enq_ready),
    .io_enq_valid(qb_q_io_enq_valid),
    .io_enq_bits_data(qb_q_io_enq_bits_data),
    .io_enq_bits_last(qb_q_io_enq_bits_last),
    .io_enq_bits_beats(qb_q_io_enq_bits_beats),
    .io_deq_ready(qb_q_io_deq_ready),
    .io_deq_valid(qb_q_io_deq_valid),
    .io_deq_bits_data(qb_q_io_deq_bits_data),
    .io_deq_bits_last(qb_q_io_deq_bits_last),
    .io_deq_bits_beats(qb_q_io_deq_bits_beats)
  );
  ShiftQueue qc_q ( // @[ShiftQueue.scala 60:19]
    .clock(qc_q_clock),
    .reset(qc_q_reset),
    .io_enq_ready(qc_q_io_enq_ready),
    .io_enq_valid(qc_q_io_enq_valid),
    .io_enq_bits_data(qc_q_io_enq_bits_data),
    .io_enq_bits_last(qc_q_io_enq_bits_last),
    .io_enq_bits_beats(qc_q_io_enq_bits_beats),
    .io_deq_ready(qc_q_io_deq_ready),
    .io_deq_valid(qc_q_io_deq_valid),
    .io_deq_bits_data(qc_q_io_deq_bits_data),
    .io_deq_bits_last(qc_q_io_deq_bits_last),
    .io_deq_bits_beats(qc_q_io_deq_bits_beats)
  );
  ShiftQueue qd_q ( // @[ShiftQueue.scala 60:19]
    .clock(qd_q_clock),
    .reset(qd_q_reset),
    .io_enq_ready(qd_q_io_enq_ready),
    .io_enq_valid(qd_q_io_enq_valid),
    .io_enq_bits_data(qd_q_io_enq_bits_data),
    .io_enq_bits_last(qd_q_io_enq_bits_last),
    .io_enq_bits_beats(qd_q_io_enq_bits_beats),
    .io_deq_ready(qd_q_io_deq_ready),
    .io_deq_valid(qd_q_io_deq_valid),
    .io_deq_bits_data(qd_q_io_deq_bits_data),
    .io_deq_bits_last(qd_q_io_deq_bits_last),
    .io_deq_bits_beats(qd_q_io_deq_bits_beats)
  );
  ShiftQueue qe_q ( // @[ShiftQueue.scala 60:19]
    .clock(qe_q_clock),
    .reset(qe_q_reset),
    .io_enq_ready(qe_q_io_enq_ready),
    .io_enq_valid(qe_q_io_enq_valid),
    .io_enq_bits_data(qe_q_io_enq_bits_data),
    .io_enq_bits_last(qe_q_io_enq_bits_last),
    .io_enq_bits_beats(qe_q_io_enq_bits_beats),
    .io_deq_ready(qe_q_io_deq_ready),
    .io_deq_valid(qe_q_io_deq_valid),
    .io_deq_bits_data(qe_q_io_deq_bits_data),
    .io_deq_bits_last(qe_q_io_deq_bits_last),
    .io_deq_bits_beats(qe_q_io_deq_bits_beats)
  );
  ShiftQueue ioX_cq ( // @[TX.scala 56:20]
    .clock(ioX_cq_clock),
    .reset(ioX_cq_reset),
    .io_enq_ready(ioX_cq_io_enq_ready),
    .io_enq_valid(ioX_cq_io_enq_valid),
    .io_enq_bits_data(ioX_cq_io_enq_bits_data),
    .io_enq_bits_last(ioX_cq_io_enq_bits_last),
    .io_enq_bits_beats(ioX_cq_io_enq_bits_beats),
    .io_deq_ready(ioX_cq_io_deq_ready),
    .io_deq_valid(ioX_cq_io_deq_valid),
    .io_deq_bits_data(ioX_cq_io_deq_bits_data),
    .io_deq_bits_last(ioX_cq_io_deq_bits_last),
    .io_deq_bits_beats(ioX_cq_io_deq_bits_beats)
  );
  ShiftQueue ioX_cq_1 ( // @[TX.scala 56:20]
    .clock(ioX_cq_1_clock),
    .reset(ioX_cq_1_reset),
    .io_enq_ready(ioX_cq_1_io_enq_ready),
    .io_enq_valid(ioX_cq_1_io_enq_valid),
    .io_enq_bits_data(ioX_cq_1_io_enq_bits_data),
    .io_enq_bits_last(ioX_cq_1_io_enq_bits_last),
    .io_enq_bits_beats(ioX_cq_1_io_enq_bits_beats),
    .io_deq_ready(ioX_cq_1_io_deq_ready),
    .io_deq_valid(ioX_cq_1_io_deq_valid),
    .io_deq_bits_data(ioX_cq_1_io_deq_bits_data),
    .io_deq_bits_last(ioX_cq_1_io_deq_bits_last),
    .io_deq_bits_beats(ioX_cq_1_io_deq_bits_beats)
  );
  ShiftQueue ioX_cq_2 ( // @[TX.scala 56:20]
    .clock(ioX_cq_2_clock),
    .reset(ioX_cq_2_reset),
    .io_enq_ready(ioX_cq_2_io_enq_ready),
    .io_enq_valid(ioX_cq_2_io_enq_valid),
    .io_enq_bits_data(ioX_cq_2_io_enq_bits_data),
    .io_enq_bits_last(ioX_cq_2_io_enq_bits_last),
    .io_enq_bits_beats(ioX_cq_2_io_enq_bits_beats),
    .io_deq_ready(ioX_cq_2_io_deq_ready),
    .io_deq_valid(ioX_cq_2_io_deq_valid),
    .io_deq_bits_data(ioX_cq_2_io_deq_bits_data),
    .io_deq_bits_last(ioX_cq_2_io_deq_bits_last),
    .io_deq_bits_beats(ioX_cq_2_io_deq_bits_beats)
  );
  ShiftQueue ioX_cq_3 ( // @[TX.scala 56:20]
    .clock(ioX_cq_3_clock),
    .reset(ioX_cq_3_reset),
    .io_enq_ready(ioX_cq_3_io_enq_ready),
    .io_enq_valid(ioX_cq_3_io_enq_valid),
    .io_enq_bits_data(ioX_cq_3_io_enq_bits_data),
    .io_enq_bits_last(ioX_cq_3_io_enq_bits_last),
    .io_enq_bits_beats(ioX_cq_3_io_enq_bits_beats),
    .io_deq_ready(ioX_cq_3_io_deq_ready),
    .io_deq_valid(ioX_cq_3_io_deq_valid),
    .io_deq_bits_data(ioX_cq_3_io_deq_bits_data),
    .io_deq_bits_last(ioX_cq_3_io_deq_bits_last),
    .io_deq_bits_beats(ioX_cq_3_io_deq_bits_beats)
  );
  ShiftQueue ioX_cq_4 ( // @[TX.scala 56:20]
    .clock(ioX_cq_4_clock),
    .reset(ioX_cq_4_reset),
    .io_enq_ready(ioX_cq_4_io_enq_ready),
    .io_enq_valid(ioX_cq_4_io_enq_valid),
    .io_enq_bits_data(ioX_cq_4_io_enq_bits_data),
    .io_enq_bits_last(ioX_cq_4_io_enq_bits_last),
    .io_enq_bits_beats(ioX_cq_4_io_enq_bits_beats),
    .io_deq_ready(ioX_cq_4_io_deq_ready),
    .io_deq_valid(ioX_cq_4_io_deq_valid),
    .io_deq_bits_data(ioX_cq_4_io_deq_bits_data),
    .io_deq_bits_last(ioX_cq_4_io_deq_bits_last),
    .io_deq_bits_beats(ioX_cq_4_io_deq_bits_beats)
  );
  ShiftQueue rxQ ( // @[TX.scala 64:19]
    .clock(rxQ_clock),
    .reset(rxQ_reset),
    .io_enq_ready(rxQ_io_enq_ready),
    .io_enq_valid(rxQ_io_enq_valid),
    .io_enq_bits_data(rxQ_io_enq_bits_data),
    .io_enq_bits_last(rxQ_io_enq_bits_last),
    .io_enq_bits_beats(rxQ_io_enq_bits_beats),
    .io_deq_ready(rxQ_io_deq_ready),
    .io_deq_valid(rxQ_io_deq_valid),
    .io_deq_bits_data(rxQ_io_deq_bits_data),
    .io_deq_bits_last(rxQ_io_deq_bits_last),
    .io_deq_bits_beats(rxQ_io_deq_bits_beats)
  );
  AsyncResetReg io_c2b_rst_reg ( // @[AsyncResetReg.scala 74:21]
    .io_q(io_c2b_rst_reg_io_q),
    .io_clk(io_c2b_rst_reg_io_clk),
    .io_rst(io_c2b_rst_reg_io_rst)
  );
  assign io_c2b_clk = clock; // @[TX.scala 122:15]
  assign io_c2b_rst = io_c2b_rst_reg_io_q; // @[TX.scala 123:15]
  assign io_c2b_send = io_c2b_send_REG_1; // @[TX.scala 124:15]
  assign io_c2b_data = io_c2b_data_REG_1; // @[TX.scala 125:15]
  assign io_sa_ready = qa_q_io_enq_ready; // @[ShiftQueue.scala 61:14]
  assign io_sb_ready = qb_q_io_enq_ready; // @[ShiftQueue.scala 61:14]
  assign io_sc_ready = qc_q_io_enq_ready; // @[ShiftQueue.scala 61:14]
  assign io_sd_ready = qd_q_io_enq_ready; // @[ShiftQueue.scala 61:14]
  assign io_rxc_ridx = rxInc_sink_io_async_ridx; // @[AsyncQueue.scala 208:19]
  assign io_rxc_safe_ridx_valid = rxInc_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 208:19]
  assign io_rxc_safe_sink_reset_n = rxInc_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 208:19]
  assign io_txc_ridx = txInc_sink_io_async_ridx; // @[AsyncQueue.scala 208:19]
  assign io_txc_safe_ridx_valid = txInc_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 208:19]
  assign io_txc_safe_sink_reset_n = txInc_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 208:19]
  assign rxInc_sink_clock = clock;
  assign rxInc_sink_reset = reset;
  assign rxInc_sink_io_deq_ready = 1'h1; // @[TX.scala 37:15]
  assign rxInc_sink_io_async_mem_0_a = io_rxc_mem_0_a; // @[AsyncQueue.scala 208:19]
  assign rxInc_sink_io_async_mem_0_b = io_rxc_mem_0_b; // @[AsyncQueue.scala 208:19]
  assign rxInc_sink_io_async_mem_0_c = io_rxc_mem_0_c; // @[AsyncQueue.scala 208:19]
  assign rxInc_sink_io_async_mem_0_d = io_rxc_mem_0_d; // @[AsyncQueue.scala 208:19]
  assign rxInc_sink_io_async_mem_0_e = io_rxc_mem_0_e; // @[AsyncQueue.scala 208:19]
  assign rxInc_sink_io_async_widx = io_rxc_widx; // @[AsyncQueue.scala 208:19]
  assign rxInc_sink_io_async_safe_widx_valid = io_rxc_safe_widx_valid; // @[AsyncQueue.scala 208:19]
  assign rxInc_sink_io_async_safe_source_reset_n = io_rxc_safe_source_reset_n; // @[AsyncQueue.scala 208:19]
  assign txInc_sink_clock = clock;
  assign txInc_sink_reset = reset;
  assign txInc_sink_io_deq_ready = 1'h1; // @[TX.scala 38:15]
  assign txInc_sink_io_async_mem_0_a = io_txc_mem_0_a; // @[AsyncQueue.scala 208:19]
  assign txInc_sink_io_async_mem_0_b = io_txc_mem_0_b; // @[AsyncQueue.scala 208:19]
  assign txInc_sink_io_async_mem_0_c = io_txc_mem_0_c; // @[AsyncQueue.scala 208:19]
  assign txInc_sink_io_async_mem_0_d = io_txc_mem_0_d; // @[AsyncQueue.scala 208:19]
  assign txInc_sink_io_async_mem_0_e = io_txc_mem_0_e; // @[AsyncQueue.scala 208:19]
  assign txInc_sink_io_async_widx = io_txc_widx; // @[AsyncQueue.scala 208:19]
  assign txInc_sink_io_async_safe_widx_valid = io_txc_safe_widx_valid; // @[AsyncQueue.scala 208:19]
  assign txInc_sink_io_async_safe_source_reset_n = io_txc_safe_source_reset_n; // @[AsyncQueue.scala 208:19]
  assign qa_q_clock = clock;
  assign qa_q_reset = reset;
  assign qa_q_io_enq_valid = io_sa_valid; // @[ShiftQueue.scala 61:14]
  assign qa_q_io_enq_bits_data = io_sa_bits_data; // @[ShiftQueue.scala 61:14]
  assign qa_q_io_enq_bits_last = io_sa_bits_last; // @[ShiftQueue.scala 61:14]
  assign qa_q_io_enq_bits_beats = io_sa_bits_beats; // @[ShiftQueue.scala 61:14]
  assign qa_q_io_deq_ready = ioX_cq_io_enq_ready & ioX_allow; // @[TX.scala 59:32]
  assign qb_q_clock = clock;
  assign qb_q_reset = reset;
  assign qb_q_io_enq_valid = 1'h0; // @[ShiftQueue.scala 61:14]
  assign qb_q_io_enq_bits_data = io_sb_bits_data; // @[ShiftQueue.scala 61:14]
  assign qb_q_io_enq_bits_last = io_sb_bits_last; // @[ShiftQueue.scala 61:14]
  assign qb_q_io_enq_bits_beats = 7'h3; // @[ShiftQueue.scala 61:14]
  assign qb_q_io_deq_ready = ioX_cq_1_io_enq_ready & ioX_allow_1; // @[TX.scala 59:32]
  assign qc_q_clock = clock;
  assign qc_q_reset = reset;
  assign qc_q_io_enq_valid = 1'h0; // @[ShiftQueue.scala 61:14]
  assign qc_q_io_enq_bits_data = io_sc_bits_data; // @[ShiftQueue.scala 61:14]
  assign qc_q_io_enq_bits_last = io_sc_bits_last; // @[ShiftQueue.scala 61:14]
  assign qc_q_io_enq_bits_beats = 7'h3; // @[ShiftQueue.scala 61:14]
  assign qc_q_io_deq_ready = ioX_cq_2_io_enq_ready & ioX_allow_2; // @[TX.scala 59:32]
  assign qd_q_clock = clock;
  assign qd_q_reset = reset;
  assign qd_q_io_enq_valid = io_sd_valid; // @[ShiftQueue.scala 61:14]
  assign qd_q_io_enq_bits_data = io_sd_bits_data; // @[ShiftQueue.scala 61:14]
  assign qd_q_io_enq_bits_last = io_sd_bits_last; // @[ShiftQueue.scala 61:14]
  assign qd_q_io_enq_bits_beats = io_sd_bits_beats; // @[ShiftQueue.scala 61:14]
  assign qd_q_io_deq_ready = ioX_cq_3_io_enq_ready & ioX_allow_3; // @[TX.scala 59:32]
  assign qe_q_clock = clock;
  assign qe_q_reset = reset;
  assign qe_q_io_enq_valid = 1'h0; // @[ShiftQueue.scala 61:14]
  assign qe_q_io_enq_bits_data = io_se_bits_data; // @[ShiftQueue.scala 61:14]
  assign qe_q_io_enq_bits_last = 1'h1; // @[ShiftQueue.scala 61:14]
  assign qe_q_io_enq_bits_beats = 7'h1; // @[ShiftQueue.scala 61:14]
  assign qe_q_io_deq_ready = ioX_cq_4_io_enq_ready & ioX_allow_4; // @[TX.scala 59:32]
  assign ioX_cq_clock = clock;
  assign ioX_cq_reset = reset;
  assign ioX_cq_io_enq_valid = qa_q_io_deq_valid & ioX_allow; // @[TX.scala 58:32]
  assign ioX_cq_io_enq_bits_data = qa_q_io_deq_bits_data; // @[TX.scala 57:20]
  assign ioX_cq_io_enq_bits_last = qa_q_io_deq_bits_last; // @[TX.scala 57:20]
  assign ioX_cq_io_enq_bits_beats = qa_q_io_deq_bits_beats; // @[TX.scala 57:20]
  assign ioX_cq_io_deq_ready = allowed[0] & ~txBusy; // @[TX.scala 100:77]
  assign ioX_cq_1_clock = clock;
  assign ioX_cq_1_reset = reset;
  assign ioX_cq_1_io_enq_valid = qb_q_io_deq_valid & ioX_allow_1; // @[TX.scala 58:32]
  assign ioX_cq_1_io_enq_bits_data = qb_q_io_deq_bits_data; // @[TX.scala 57:20]
  assign ioX_cq_1_io_enq_bits_last = qb_q_io_deq_bits_last; // @[TX.scala 57:20]
  assign ioX_cq_1_io_enq_bits_beats = qb_q_io_deq_bits_beats; // @[TX.scala 57:20]
  assign ioX_cq_1_io_deq_ready = allowed[1] & ~txBusy; // @[TX.scala 100:77]
  assign ioX_cq_2_clock = clock;
  assign ioX_cq_2_reset = reset;
  assign ioX_cq_2_io_enq_valid = qc_q_io_deq_valid & ioX_allow_2; // @[TX.scala 58:32]
  assign ioX_cq_2_io_enq_bits_data = qc_q_io_deq_bits_data; // @[TX.scala 57:20]
  assign ioX_cq_2_io_enq_bits_last = qc_q_io_deq_bits_last; // @[TX.scala 57:20]
  assign ioX_cq_2_io_enq_bits_beats = qc_q_io_deq_bits_beats; // @[TX.scala 57:20]
  assign ioX_cq_2_io_deq_ready = allowed[2] & ~txBusy; // @[TX.scala 100:77]
  assign ioX_cq_3_clock = clock;
  assign ioX_cq_3_reset = reset;
  assign ioX_cq_3_io_enq_valid = qd_q_io_deq_valid & ioX_allow_3; // @[TX.scala 58:32]
  assign ioX_cq_3_io_enq_bits_data = qd_q_io_deq_bits_data; // @[TX.scala 57:20]
  assign ioX_cq_3_io_enq_bits_last = qd_q_io_deq_bits_last; // @[TX.scala 57:20]
  assign ioX_cq_3_io_enq_bits_beats = qd_q_io_deq_bits_beats; // @[TX.scala 57:20]
  assign ioX_cq_3_io_deq_ready = allowed[3] & ~txBusy; // @[TX.scala 100:77]
  assign ioX_cq_4_clock = clock;
  assign ioX_cq_4_reset = reset;
  assign ioX_cq_4_io_enq_valid = qe_q_io_deq_valid & ioX_allow_4; // @[TX.scala 58:32]
  assign ioX_cq_4_io_enq_bits_data = qe_q_io_deq_bits_data; // @[TX.scala 57:20]
  assign ioX_cq_4_io_enq_bits_last = qe_q_io_deq_bits_last; // @[TX.scala 57:20]
  assign ioX_cq_4_io_enq_bits_beats = qe_q_io_deq_bits_beats; // @[TX.scala 57:20]
  assign ioX_cq_4_io_deq_ready = allowed[4] & ~txBusy; // @[TX.scala 100:77]
  assign rxQ_clock = clock;
  assign rxQ_reset = reset;
  assign rxQ_io_enq_valid = |rxHeader[31:7]; // @[TX.scala 66:42]
  assign rxQ_io_enq_bits_data = {header_hi,header_lo}; // @[Cat.scala 30:58]
  assign rxQ_io_enq_bits_last = 1'h1; // @[TX.scala 68:25]
  assign rxQ_io_enq_bits_beats = 7'h1; // @[TX.scala 69:25]
  assign rxQ_io_deq_ready = f_ready & allowReturn; // @[TX.scala 89:31]
  assign io_c2b_rst_reg_io_clk = clock; // @[AsyncResetReg.scala 76:16]
  assign io_c2b_rst_reg_io_rst = reset; // @[compatibility.scala 260:56]
  always @(posedge clock) begin
    if (reset) begin // @[TX.scala 31:19]
      rx_a <= 20'h0; // @[TX.scala 31:19]
    end else begin
      rx_a <= rx_out_2_a; // @[TX.scala 70:6]
    end
    if (reset) begin // @[TX.scala 31:19]
      rx_b <= 20'h0; // @[TX.scala 31:19]
    end else begin
      rx_b <= rx_out_2_b; // @[TX.scala 70:6]
    end
    if (reset) begin // @[TX.scala 31:19]
      rx_c <= 20'h0; // @[TX.scala 31:19]
    end else begin
      rx_c <= rx_out_2_c; // @[TX.scala 70:6]
    end
    if (reset) begin // @[TX.scala 31:19]
      rx_d <= 20'h0; // @[TX.scala 31:19]
    end else begin
      rx_d <= rx_out_2_d; // @[TX.scala 70:6]
    end
    if (reset) begin // @[TX.scala 31:19]
      rx_e <= 20'h0; // @[TX.scala 31:19]
    end else begin
      rx_e <= rx_out_2_e; // @[TX.scala 70:6]
    end
    if (reset) begin // @[TX.scala 32:19]
      tx_a <= 20'h0; // @[TX.scala 32:19]
    end else begin
      tx_a <= _ioX_tx_a_T_6[19:0]; // @[TX.scala 54:12]
    end
    if (reset) begin // @[TX.scala 32:19]
      tx_b <= 20'h0; // @[TX.scala 32:19]
    end else begin
      tx_b <= _ioX_tx_bT_6[19:0]; // @[TX.scala 54:12]
    end
    if (reset) begin // @[TX.scala 32:19]
      tx_c <= 20'h0; // @[TX.scala 32:19]
    end else begin
      tx_c <= _ioX_tx_c_T_6[19:0]; // @[TX.scala 54:12]
    end
    if (reset) begin // @[TX.scala 32:19]
      tx_d <= 20'h0; // @[TX.scala 32:19]
    end else begin
      tx_d <= _ioX_tx_d_T_6[19:0]; // @[TX.scala 54:12]
    end
    if (reset) begin // @[TX.scala 32:19]
      tx_e <= 20'h0; // @[TX.scala 32:19]
    end else begin
      tx_e <= _ioX_tx_e_T_6[19:0]; // @[TX.scala 54:12]
    end
    ioX_first <= reset | _GEN_0; // @[Reg.scala 27:20 Reg.scala 27:20]
    ioX_first_1 <= reset | _GEN_1; // @[Reg.scala 27:20 Reg.scala 27:20]
    ioX_first_2 <= reset | _GEN_2; // @[Reg.scala 27:20 Reg.scala 27:20]
    ioX_first_3 <= reset | _GEN_3; // @[Reg.scala 27:20 Reg.scala 27:20]
    ioX_first_4 <= reset | _GEN_4; // @[Reg.scala 27:20 Reg.scala 27:20]
    if (reset) begin // @[TX.scala 80:21]
      xmit <= 2'h0; // @[TX.scala 80:21]
    end else if (_T_1) begin // @[TX.scala 83:19]
      xmit <= 2'h3; // @[TX.scala 83:26]
    end else if (~forceXmit) begin // @[TX.scala 82:21]
      xmit <= _xmit_T_1; // @[TX.scala 82:28]
    end
    first <= reset | _GEN_8; // @[TX.scala 92:22 TX.scala 92:22]
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask <= 6'h3f; // @[Arbiter.scala 23:23]
    end else if (first & |requests) begin // @[Arbiter.scala 27:32]
      readys_mask <= _readys_mask_T_9; // @[Arbiter.scala 28:12]
    end
    if (first) begin // @[TX.scala 106:16]
      state <= _readys_mask_T; // @[TX.scala 106:24]
    end
    if (reset) begin // @[TX.scala 99:23]
      txBusy <= 1'h0; // @[TX.scala 99:23]
    end else if (txBusy) begin // @[TX.scala 112:16]
      if (transferByteCnt == 2'h3) begin // @[TX.scala 114:35]
        txBusy <= 1'h0; // @[TX.scala 115:14]
      end else begin
        txBusy <= _GEN_10;
      end
    end else begin
      txBusy <= _GEN_10;
    end
    if (reset) begin // @[TX.scala 108:32]
      transferByteCnt <= 2'h0; // @[TX.scala 108:32]
    end else if (txBusy) begin // @[TX.scala 112:16]
      transferByteCnt <= _transferByteCnt_T_1; // @[TX.scala 113:21]
    end
    if (send) begin // @[Reg.scala 16:19]
      transferDataReg <= _transferDataReg_T_16; // @[Reg.scala 16:23]
    end
    io_c2b_send_REG <= txBusy; // @[TX.scala 124:33]
    io_c2b_send_REG_1 <= io_c2b_send_REG; // @[TX.scala 124:25]
    if (2'h3 == transferByteCnt) begin // @[TX.scala 125:33]
      io_c2b_data_REG <= transferBytes_3; // @[TX.scala 125:33]
    end else if (2'h2 == transferByteCnt) begin // @[TX.scala 125:33]
      io_c2b_data_REG <= transferBytes_2; // @[TX.scala 125:33]
    end else if (2'h1 == transferByteCnt) begin // @[TX.scala 125:33]
      io_c2b_data_REG <= transferBytes_1; // @[TX.scala 125:33]
    end else begin
      io_c2b_data_REG <= transferBytes_0;
    end
    io_c2b_data_REG_1 <= io_c2b_data_REG; // @[TX.scala 125:25]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rx_a = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  rx_b = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  rx_c = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  rx_d = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  rx_e = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  tx_a = _RAND_5[19:0];
  _RAND_6 = {1{`RANDOM}};
  tx_b = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  tx_c = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  tx_d = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  tx_e = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  ioX_first = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ioX_first_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ioX_first_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ioX_first_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ioX_first_4 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  xmit = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  first = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  readys_mask = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  state = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  txBusy = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  transferByteCnt = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  transferDataReg = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  io_c2b_send_REG = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  io_c2b_send_REG_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  io_c2b_data_REG = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  io_c2b_data_REG_1 = _RAND_25[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ResetCatchAndSync_d3(
  input   clock,
  input   reset,
  output  io_sync_reset
);
  wire  io_sync_reset_chain_clock; // @[ShiftReg.scala 45:23]
  wire  io_sync_reset_chain_reset; // @[ShiftReg.scala 45:23]
  wire  io_sync_reset_chain_io_d; // @[ShiftReg.scala 45:23]
  wire  io_sync_reset_chain_io_q; // @[ShiftReg.scala 45:23]
  wire  _io_sync_reset_WIRE = io_sync_reset_chain_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  AsyncResetSynchronizerShiftReg_w1_d3_i0_20 io_sync_reset_chain ( // @[ShiftReg.scala 45:23]
    .clock(io_sync_reset_chain_clock),
    .reset(io_sync_reset_chain_reset),
    .io_d(io_sync_reset_chain_io_d),
    .io_q(io_sync_reset_chain_io_q)
  );
  assign io_sync_reset = ~_io_sync_reset_WIRE; // @[ResetCatchAndSync.scala 29:7]
  assign io_sync_reset_chain_clock = clock;
  assign io_sync_reset_chain_reset = reset; // @[ResetCatchAndSync.scala 26:27]
  assign io_sync_reset_chain_io_d = 1'h1; // @[ShiftReg.scala 47:16]
endmodule
module ChipLink(
  input         clock,
  input         reset,
  input         auto_mbypass_out_a_ready,
  output        auto_mbypass_out_a_valid,
  output [2:0]  auto_mbypass_out_a_bits_opcode,
  output [2:0]  auto_mbypass_out_a_bits_param,
  output [2:0]  auto_mbypass_out_a_bits_size,
  output [5:0]  auto_mbypass_out_a_bits_source,
  output [31:0] auto_mbypass_out_a_bits_address,
  output [3:0]  auto_mbypass_out_a_bits_mask,
  output [31:0] auto_mbypass_out_a_bits_data,
  input         auto_mbypass_out_c_ready,
  output        auto_mbypass_out_c_valid,
  output [2:0]  auto_mbypass_out_c_bits_opcode,
  output [2:0]  auto_mbypass_out_c_bits_param,
  output [2:0]  auto_mbypass_out_c_bits_size,
  output [5:0]  auto_mbypass_out_c_bits_source,
  output [31:0] auto_mbypass_out_c_bits_address,
  output        auto_mbypass_out_d_ready,
  input         auto_mbypass_out_d_valid,
  input  [2:0]  auto_mbypass_out_d_bits_opcode,
  input  [1:0]  auto_mbypass_out_d_bits_param,
  input  [2:0]  auto_mbypass_out_d_bits_size,
  input  [5:0]  auto_mbypass_out_d_bits_source,
  input         auto_mbypass_out_d_bits_denied,
  input  [31:0] auto_mbypass_out_d_bits_data,
  input         auto_mbypass_out_d_bits_corrupt,
  input         auto_mbypass_out_e_ready,
  output        auto_mbypass_out_e_valid,
  output        auto_mbypass_out_e_bits_sink,
  output        auto_sbypass_node_in_in_a_ready,
  input         auto_sbypass_node_in_in_a_valid,
  input  [2:0]  auto_sbypass_node_in_in_a_bits_opcode,
  input  [2:0]  auto_sbypass_node_in_in_a_bits_size,
  input  [3:0]  auto_sbypass_node_in_in_a_bits_source,
  input  [31:0] auto_sbypass_node_in_in_a_bits_address,
  input  [3:0]  auto_sbypass_node_in_in_a_bits_mask,
  input  [31:0] auto_sbypass_node_in_in_a_bits_data,
  input         auto_sbypass_node_in_in_d_ready,
  output        auto_sbypass_node_in_in_d_valid,
  output [2:0]  auto_sbypass_node_in_in_d_bits_opcode,
  output [1:0]  auto_sbypass_node_in_in_d_bits_param,
  output [2:0]  auto_sbypass_node_in_in_d_bits_size,
  output [3:0]  auto_sbypass_node_in_in_d_bits_source,
  output [4:0]  auto_sbypass_node_in_in_d_bits_sink,
  output        auto_sbypass_node_in_in_d_bits_denied,
  output [31:0] auto_sbypass_node_in_in_d_bits_data,
  output        auto_sbypass_node_in_in_d_bits_corrupt,
  output        auto_io_out_c2b_clk,
  output        auto_io_out_c2b_rst,
  output        auto_io_out_c2b_send,
  output [7:0]  auto_io_out_c2b_data,
  input         auto_io_out_b2c_clk,
  input         auto_io_out_b2c_rst,
  input         auto_io_out_b2c_send,
  input  [7:0]  auto_io_out_b2c_data
);
  wire  sbypass_clock; // @[ChipLink.scala 65:35]
  wire  sbypass_reset; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_out_out_a_ready; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_out_out_a_valid; // @[ChipLink.scala 65:35]
  wire [2:0] sbypass_auto_node_out_out_a_bits_opcode; // @[ChipLink.scala 65:35]
  wire [2:0] sbypass_auto_node_out_out_a_bits_size; // @[ChipLink.scala 65:35]
  wire [3:0] sbypass_auto_node_out_out_a_bits_source; // @[ChipLink.scala 65:35]
  wire [31:0] sbypass_auto_node_out_out_a_bits_address; // @[ChipLink.scala 65:35]
  wire [3:0] sbypass_auto_node_out_out_a_bits_mask; // @[ChipLink.scala 65:35]
  wire [31:0] sbypass_auto_node_out_out_a_bits_data; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_out_out_d_ready; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_out_out_d_valid; // @[ChipLink.scala 65:35]
  wire [2:0] sbypass_auto_node_out_out_d_bits_opcode; // @[ChipLink.scala 65:35]
  wire [1:0] sbypass_auto_node_out_out_d_bits_param; // @[ChipLink.scala 65:35]
  wire [2:0] sbypass_auto_node_out_out_d_bits_size; // @[ChipLink.scala 65:35]
  wire [3:0] sbypass_auto_node_out_out_d_bits_source; // @[ChipLink.scala 65:35]
  wire [4:0] sbypass_auto_node_out_out_d_bits_sink; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_out_out_d_bits_denied; // @[ChipLink.scala 65:35]
  wire [31:0] sbypass_auto_node_out_out_d_bits_data; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_out_out_d_bits_corrupt; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_in_in_a_ready; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_in_in_a_valid; // @[ChipLink.scala 65:35]
  wire [2:0] sbypass_auto_node_in_in_a_bits_opcode; // @[ChipLink.scala 65:35]
  wire [2:0] sbypass_auto_node_in_in_a_bits_size; // @[ChipLink.scala 65:35]
  wire [3:0] sbypass_auto_node_in_in_a_bits_source; // @[ChipLink.scala 65:35]
  wire [31:0] sbypass_auto_node_in_in_a_bits_address; // @[ChipLink.scala 65:35]
  wire [3:0] sbypass_auto_node_in_in_a_bits_mask; // @[ChipLink.scala 65:35]
  wire [31:0] sbypass_auto_node_in_in_a_bits_data; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_in_in_d_ready; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_in_in_d_valid; // @[ChipLink.scala 65:35]
  wire [2:0] sbypass_auto_node_in_in_d_bits_opcode; // @[ChipLink.scala 65:35]
  wire [1:0] sbypass_auto_node_in_in_d_bits_param; // @[ChipLink.scala 65:35]
  wire [2:0] sbypass_auto_node_in_in_d_bits_size; // @[ChipLink.scala 65:35]
  wire [3:0] sbypass_auto_node_in_in_d_bits_source; // @[ChipLink.scala 65:35]
  wire [4:0] sbypass_auto_node_in_in_d_bits_sink; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_in_in_d_bits_denied; // @[ChipLink.scala 65:35]
  wire [31:0] sbypass_auto_node_in_in_d_bits_data; // @[ChipLink.scala 65:35]
  wire  sbypass_auto_node_in_in_d_bits_corrupt; // @[ChipLink.scala 65:35]
  wire  sbypass_io_bypass; // @[ChipLink.scala 65:35]
  wire  mbypass_clock; // @[ChipLink.scala 69:35]
  wire  mbypass_reset; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_a_ready; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_a_valid; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_in_1_a_bits_opcode; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_in_1_a_bits_param; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_in_1_a_bits_size; // @[ChipLink.scala 69:35]
  wire [5:0] mbypass_auto_in_1_a_bits_source; // @[ChipLink.scala 69:35]
  wire [31:0] mbypass_auto_in_1_a_bits_address; // @[ChipLink.scala 69:35]
  wire [3:0] mbypass_auto_in_1_a_bits_mask; // @[ChipLink.scala 69:35]
  wire [31:0] mbypass_auto_in_1_a_bits_data; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_c_ready; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_c_valid; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_in_1_c_bits_opcode; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_in_1_c_bits_param; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_in_1_c_bits_size; // @[ChipLink.scala 69:35]
  wire [5:0] mbypass_auto_in_1_c_bits_source; // @[ChipLink.scala 69:35]
  wire [31:0] mbypass_auto_in_1_c_bits_address; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_d_ready; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_d_valid; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_in_1_d_bits_opcode; // @[ChipLink.scala 69:35]
  wire [1:0] mbypass_auto_in_1_d_bits_param; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_in_1_d_bits_size; // @[ChipLink.scala 69:35]
  wire [5:0] mbypass_auto_in_1_d_bits_source; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_d_bits_denied; // @[ChipLink.scala 69:35]
  wire [31:0] mbypass_auto_in_1_d_bits_data; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_e_ready; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_e_valid; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_in_1_e_bits_sink; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_a_ready; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_a_valid; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_out_a_bits_opcode; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_out_a_bits_param; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_out_a_bits_size; // @[ChipLink.scala 69:35]
  wire [5:0] mbypass_auto_out_a_bits_source; // @[ChipLink.scala 69:35]
  wire [31:0] mbypass_auto_out_a_bits_address; // @[ChipLink.scala 69:35]
  wire [3:0] mbypass_auto_out_a_bits_mask; // @[ChipLink.scala 69:35]
  wire [31:0] mbypass_auto_out_a_bits_data; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_c_ready; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_c_valid; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_out_c_bits_opcode; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_out_c_bits_param; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_out_c_bits_size; // @[ChipLink.scala 69:35]
  wire [5:0] mbypass_auto_out_c_bits_source; // @[ChipLink.scala 69:35]
  wire [31:0] mbypass_auto_out_c_bits_address; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_d_ready; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_d_valid; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_out_d_bits_opcode; // @[ChipLink.scala 69:35]
  wire [1:0] mbypass_auto_out_d_bits_param; // @[ChipLink.scala 69:35]
  wire [2:0] mbypass_auto_out_d_bits_size; // @[ChipLink.scala 69:35]
  wire [5:0] mbypass_auto_out_d_bits_source; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_d_bits_denied; // @[ChipLink.scala 69:35]
  wire [31:0] mbypass_auto_out_d_bits_data; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_d_bits_corrupt; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_e_ready; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_e_valid; // @[ChipLink.scala 69:35]
  wire  mbypass_auto_out_e_bits_sink; // @[ChipLink.scala 69:35]
  wire  mbypass_io_bypass; // @[ChipLink.scala 69:35]
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire [4:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  sinkA_clock; // @[ChipLink.scala 148:23]
  wire  sinkA_reset; // @[ChipLink.scala 148:23]
  wire  sinkA_io_a_ready; // @[ChipLink.scala 148:23]
  wire  sinkA_io_a_valid; // @[ChipLink.scala 148:23]
  wire [2:0] sinkA_io_a_bits_opcode; // @[ChipLink.scala 148:23]
  wire [2:0] sinkA_io_a_bits_size; // @[ChipLink.scala 148:23]
  wire [3:0] sinkA_io_a_bits_source; // @[ChipLink.scala 148:23]
  wire [31:0] sinkA_io_a_bits_address; // @[ChipLink.scala 148:23]
  wire [3:0] sinkA_io_a_bits_mask; // @[ChipLink.scala 148:23]
  wire [31:0] sinkA_io_a_bits_data; // @[ChipLink.scala 148:23]
  wire  sinkA_io_q_ready; // @[ChipLink.scala 148:23]
  wire  sinkA_io_q_valid; // @[ChipLink.scala 148:23]
  wire [31:0] sinkA_io_q_bits_data; // @[ChipLink.scala 148:23]
  wire  sinkA_io_q_bits_last; // @[ChipLink.scala 148:23]
  wire [6:0] sinkA_io_q_bits_beats; // @[ChipLink.scala 148:23]
  wire  sinkB_clock; // @[ChipLink.scala 149:23]
  wire  sinkB_reset; // @[ChipLink.scala 149:23]
  wire  sinkB_io_q_ready; // @[ChipLink.scala 149:23]
  wire  sinkB_io_q_valid; // @[ChipLink.scala 149:23]
  wire [31:0] sinkB_io_q_bits_data; // @[ChipLink.scala 149:23]
  wire  sinkB_io_q_bits_last; // @[ChipLink.scala 149:23]
  wire  sinkC_clock; // @[ChipLink.scala 150:23]
  wire  sinkC_reset; // @[ChipLink.scala 150:23]
  wire  sinkC_io_q_ready; // @[ChipLink.scala 150:23]
  wire  sinkC_io_q_valid; // @[ChipLink.scala 150:23]
  wire [31:0] sinkC_io_q_bits_data; // @[ChipLink.scala 150:23]
  wire  sinkC_io_q_bits_last; // @[ChipLink.scala 150:23]
  wire  sinkD_clock; // @[ChipLink.scala 151:23]
  wire  sinkD_reset; // @[ChipLink.scala 151:23]
  wire  sinkD_io_d_ready; // @[ChipLink.scala 151:23]
  wire  sinkD_io_d_valid; // @[ChipLink.scala 151:23]
  wire [2:0] sinkD_io_d_bits_opcode; // @[ChipLink.scala 151:23]
  wire [1:0] sinkD_io_d_bits_param; // @[ChipLink.scala 151:23]
  wire [2:0] sinkD_io_d_bits_size; // @[ChipLink.scala 151:23]
  wire [5:0] sinkD_io_d_bits_source; // @[ChipLink.scala 151:23]
  wire  sinkD_io_d_bits_denied; // @[ChipLink.scala 151:23]
  wire [31:0] sinkD_io_d_bits_data; // @[ChipLink.scala 151:23]
  wire  sinkD_io_q_ready; // @[ChipLink.scala 151:23]
  wire  sinkD_io_q_valid; // @[ChipLink.scala 151:23]
  wire [31:0] sinkD_io_q_bits_data; // @[ChipLink.scala 151:23]
  wire  sinkD_io_q_bits_last; // @[ChipLink.scala 151:23]
  wire [6:0] sinkD_io_q_bits_beats; // @[ChipLink.scala 151:23]
  wire  sinkD_io_a_tlSource_valid; // @[ChipLink.scala 151:23]
  wire [5:0] sinkD_io_a_tlSource_bits; // @[ChipLink.scala 151:23]
  wire [15:0] sinkD_io_a_clSource; // @[ChipLink.scala 151:23]
  wire  sinkD_io_c_tlSource_valid; // @[ChipLink.scala 151:23]
  wire [5:0] sinkD_io_c_tlSource_bits; // @[ChipLink.scala 151:23]
  wire [15:0] sinkD_io_c_clSource; // @[ChipLink.scala 151:23]
  wire [31:0] sinkE_io_q_bits_data; // @[ChipLink.scala 152:23]
  wire [15:0] sinkE_io_d_clSink; // @[ChipLink.scala 152:23]
  wire  sourceA_clock; // @[ChipLink.scala 153:25]
  wire  sourceA_reset; // @[ChipLink.scala 153:25]
  wire  sourceA_io_a_ready; // @[ChipLink.scala 153:25]
  wire  sourceA_io_a_valid; // @[ChipLink.scala 153:25]
  wire [2:0] sourceA_io_a_bits_opcode; // @[ChipLink.scala 153:25]
  wire [2:0] sourceA_io_a_bits_param; // @[ChipLink.scala 153:25]
  wire [2:0] sourceA_io_a_bits_size; // @[ChipLink.scala 153:25]
  wire [5:0] sourceA_io_a_bits_source; // @[ChipLink.scala 153:25]
  wire [31:0] sourceA_io_a_bits_address; // @[ChipLink.scala 153:25]
  wire [3:0] sourceA_io_a_bits_mask; // @[ChipLink.scala 153:25]
  wire [31:0] sourceA_io_a_bits_data; // @[ChipLink.scala 153:25]
  wire  sourceA_io_q_ready; // @[ChipLink.scala 153:25]
  wire  sourceA_io_q_valid; // @[ChipLink.scala 153:25]
  wire [31:0] sourceA_io_q_bits; // @[ChipLink.scala 153:25]
  wire  sourceA_io_d_tlSource_valid; // @[ChipLink.scala 153:25]
  wire [5:0] sourceA_io_d_tlSource_bits; // @[ChipLink.scala 153:25]
  wire [15:0] sourceA_io_d_clSource; // @[ChipLink.scala 153:25]
  wire  sourceB_clock; // @[ChipLink.scala 154:25]
  wire  sourceB_reset; // @[ChipLink.scala 154:25]
  wire  sourceB_io_q_ready; // @[ChipLink.scala 154:25]
  wire  sourceB_io_q_valid; // @[ChipLink.scala 154:25]
  wire [31:0] sourceB_io_q_bits; // @[ChipLink.scala 154:25]
  wire  sourceC_clock; // @[ChipLink.scala 155:25]
  wire  sourceC_reset; // @[ChipLink.scala 155:25]
  wire  sourceC_io_c_ready; // @[ChipLink.scala 155:25]
  wire  sourceC_io_c_valid; // @[ChipLink.scala 155:25]
  wire [2:0] sourceC_io_c_bits_opcode; // @[ChipLink.scala 155:25]
  wire [2:0] sourceC_io_c_bits_param; // @[ChipLink.scala 155:25]
  wire [2:0] sourceC_io_c_bits_size; // @[ChipLink.scala 155:25]
  wire [5:0] sourceC_io_c_bits_source; // @[ChipLink.scala 155:25]
  wire [31:0] sourceC_io_c_bits_address; // @[ChipLink.scala 155:25]
  wire  sourceC_io_q_ready; // @[ChipLink.scala 155:25]
  wire  sourceC_io_q_valid; // @[ChipLink.scala 155:25]
  wire [31:0] sourceC_io_q_bits; // @[ChipLink.scala 155:25]
  wire  sourceC_io_d_tlSource_valid; // @[ChipLink.scala 155:25]
  wire [5:0] sourceC_io_d_tlSource_bits; // @[ChipLink.scala 155:25]
  wire [15:0] sourceC_io_d_clSource; // @[ChipLink.scala 155:25]
  wire  sourceD_clock; // @[ChipLink.scala 156:25]
  wire  sourceD_reset; // @[ChipLink.scala 156:25]
  wire  sourceD_io_d_ready; // @[ChipLink.scala 156:25]
  wire  sourceD_io_d_valid; // @[ChipLink.scala 156:25]
  wire [2:0] sourceD_io_d_bits_opcode; // @[ChipLink.scala 156:25]
  wire [1:0] sourceD_io_d_bits_param; // @[ChipLink.scala 156:25]
  wire [2:0] sourceD_io_d_bits_size; // @[ChipLink.scala 156:25]
  wire [3:0] sourceD_io_d_bits_source; // @[ChipLink.scala 156:25]
  wire [4:0] sourceD_io_d_bits_sink; // @[ChipLink.scala 156:25]
  wire  sourceD_io_d_bits_denied; // @[ChipLink.scala 156:25]
  wire [31:0] sourceD_io_d_bits_data; // @[ChipLink.scala 156:25]
  wire  sourceD_io_d_bits_corrupt; // @[ChipLink.scala 156:25]
  wire  sourceD_io_q_ready; // @[ChipLink.scala 156:25]
  wire  sourceD_io_q_valid; // @[ChipLink.scala 156:25]
  wire [31:0] sourceD_io_q_bits; // @[ChipLink.scala 156:25]
  wire [15:0] sourceD_io_e_clSink; // @[ChipLink.scala 156:25]
  wire  sourceE_io_e_ready; // @[ChipLink.scala 157:25]
  wire  sourceE_io_e_valid; // @[ChipLink.scala 157:25]
  wire  sourceE_io_e_bits_sink; // @[ChipLink.scala 157:25]
  wire  sourceE_io_q_ready; // @[ChipLink.scala 157:25]
  wire  sourceE_io_q_valid; // @[ChipLink.scala 157:25]
  wire [31:0] sourceE_io_q_bits; // @[ChipLink.scala 157:25]
  wire  rx_clock; // @[ChipLink.scala 159:20]
  wire  rx_reset; // @[ChipLink.scala 159:20]
  wire  rx_io_b2c_send; // @[ChipLink.scala 159:20]
  wire [7:0] rx_io_b2c_data; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_a_mem_0; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_a_mem_1; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_a_mem_2; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_a_mem_3; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_a_mem_4; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_a_mem_5; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_a_mem_6; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_a_mem_7; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_a_ridx; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_a_widx; // @[ChipLink.scala 159:20]
  wire  rx_io_a_safe_ridx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_a_safe_widx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_a_safe_source_reset_n; // @[ChipLink.scala 159:20]
  wire  rx_io_a_safe_sink_reset_n; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_bmem_0; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_bmem_1; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_bmem_2; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_bmem_3; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_bmem_4; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_bmem_5; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_bmem_6; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_bmem_7; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_bridx; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_bwidx; // @[ChipLink.scala 159:20]
  wire  rx_io_bsafe_ridx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_bsafe_widx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_bsafe_source_reset_n; // @[ChipLink.scala 159:20]
  wire  rx_io_bsafe_sink_reset_n; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_c_mem_0; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_c_mem_1; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_c_mem_2; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_c_mem_3; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_c_mem_4; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_c_mem_5; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_c_mem_6; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_c_mem_7; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_c_ridx; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_c_widx; // @[ChipLink.scala 159:20]
  wire  rx_io_c_safe_ridx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_c_safe_widx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_c_safe_source_reset_n; // @[ChipLink.scala 159:20]
  wire  rx_io_c_safe_sink_reset_n; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_d_mem_0; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_d_mem_1; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_d_mem_2; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_d_mem_3; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_d_mem_4; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_d_mem_5; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_d_mem_6; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_d_mem_7; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_d_ridx; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_d_widx; // @[ChipLink.scala 159:20]
  wire  rx_io_d_safe_ridx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_d_safe_widx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_d_safe_source_reset_n; // @[ChipLink.scala 159:20]
  wire  rx_io_d_safe_sink_reset_n; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_e_mem_0; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_e_mem_1; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_e_mem_2; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_e_mem_3; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_e_mem_4; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_e_mem_5; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_e_mem_6; // @[ChipLink.scala 159:20]
  wire [31:0] rx_io_e_mem_7; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_e_ridx; // @[ChipLink.scala 159:20]
  wire [3:0] rx_io_e_widx; // @[ChipLink.scala 159:20]
  wire  rx_io_e_safe_ridx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_e_safe_widx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_e_safe_source_reset_n; // @[ChipLink.scala 159:20]
  wire  rx_io_e_safe_sink_reset_n; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_rxc_mem_0_a; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_rxc_mem_0_b; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_rxc_mem_0_c; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_rxc_mem_0_d; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_rxc_mem_0_e; // @[ChipLink.scala 159:20]
  wire  rx_io_rxc_ridx; // @[ChipLink.scala 159:20]
  wire  rx_io_rxc_widx; // @[ChipLink.scala 159:20]
  wire  rx_io_rxc_safe_ridx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_rxc_safe_widx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_rxc_safe_source_reset_n; // @[ChipLink.scala 159:20]
  wire  rx_io_rxc_safe_sink_reset_n; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_txc_mem_0_a; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_txc_mem_0_b; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_txc_mem_0_c; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_txc_mem_0_d; // @[ChipLink.scala 159:20]
  wire [19:0] rx_io_txc_mem_0_e; // @[ChipLink.scala 159:20]
  wire  rx_io_txc_ridx; // @[ChipLink.scala 159:20]
  wire  rx_io_txc_widx; // @[ChipLink.scala 159:20]
  wire  rx_io_txc_safe_ridx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_txc_safe_widx_valid; // @[ChipLink.scala 159:20]
  wire  rx_io_txc_safe_source_reset_n; // @[ChipLink.scala 159:20]
  wire  rx_io_txc_safe_sink_reset_n; // @[ChipLink.scala 159:20]
  wire  rx_reset_reg_io_q; // @[AsyncResetReg.scala 74:21]
  wire  rx_reset_reg_io_clk; // @[AsyncResetReg.scala 74:21]
  wire  rx_reset_reg_io_rst; // @[AsyncResetReg.scala 74:21]
  wire  sourceA_io_q_sink_clock; // @[AsyncQueue.scala 207:22]
  wire  sourceA_io_q_sink_reset; // @[AsyncQueue.scala 207:22]
  wire  sourceA_io_q_sink_io_deq_ready; // @[AsyncQueue.scala 207:22]
  wire  sourceA_io_q_sink_io_deq_valid; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_deq_bits; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_async_mem_0; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_async_mem_1; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_async_mem_2; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_async_mem_3; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_async_mem_4; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_async_mem_5; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_async_mem_6; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceA_io_q_sink_io_async_mem_7; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceA_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceA_io_q_sink_io_async_widx; // @[AsyncQueue.scala 207:22]
  wire  sourceA_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceA_io_q_sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceA_io_q_sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceA_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceB_io_q_sink_clock; // @[AsyncQueue.scala 207:22]
  wire  sourceB_io_q_sink_reset; // @[AsyncQueue.scala 207:22]
  wire  sourceB_io_q_sink_io_deq_ready; // @[AsyncQueue.scala 207:22]
  wire  sourceB_io_q_sink_io_deq_valid; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_deq_bits; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_async_mem_0; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_async_mem_1; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_async_mem_2; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_async_mem_3; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_async_mem_4; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_async_mem_5; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_async_mem_6; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceB_io_q_sink_io_async_mem_7; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceB_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceB_io_q_sink_io_async_widx; // @[AsyncQueue.scala 207:22]
  wire  sourceB_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceB_io_q_sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceB_io_q_sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceB_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceC_io_q_sink_clock; // @[AsyncQueue.scala 207:22]
  wire  sourceC_io_q_sink_reset; // @[AsyncQueue.scala 207:22]
  wire  sourceC_io_q_sink_io_deq_ready; // @[AsyncQueue.scala 207:22]
  wire  sourceC_io_q_sink_io_deq_valid; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_deq_bits; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_async_mem_0; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_async_mem_1; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_async_mem_2; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_async_mem_3; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_async_mem_4; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_async_mem_5; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_async_mem_6; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceC_io_q_sink_io_async_mem_7; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceC_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceC_io_q_sink_io_async_widx; // @[AsyncQueue.scala 207:22]
  wire  sourceC_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceC_io_q_sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceC_io_q_sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceC_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceD_io_q_sink_clock; // @[AsyncQueue.scala 207:22]
  wire  sourceD_io_q_sink_reset; // @[AsyncQueue.scala 207:22]
  wire  sourceD_io_q_sink_io_deq_ready; // @[AsyncQueue.scala 207:22]
  wire  sourceD_io_q_sink_io_deq_valid; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_deq_bits; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_async_mem_0; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_async_mem_1; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_async_mem_2; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_async_mem_3; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_async_mem_4; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_async_mem_5; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_async_mem_6; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceD_io_q_sink_io_async_mem_7; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceD_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceD_io_q_sink_io_async_widx; // @[AsyncQueue.scala 207:22]
  wire  sourceD_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceD_io_q_sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceD_io_q_sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceD_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceE_io_q_sink_clock; // @[AsyncQueue.scala 207:22]
  wire  sourceE_io_q_sink_reset; // @[AsyncQueue.scala 207:22]
  wire  sourceE_io_q_sink_io_deq_ready; // @[AsyncQueue.scala 207:22]
  wire  sourceE_io_q_sink_io_deq_valid; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_deq_bits; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_async_mem_0; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_async_mem_1; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_async_mem_2; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_async_mem_3; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_async_mem_4; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_async_mem_5; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_async_mem_6; // @[AsyncQueue.scala 207:22]
  wire [31:0] sourceE_io_q_sink_io_async_mem_7; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceE_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 207:22]
  wire [3:0] sourceE_io_q_sink_io_async_widx; // @[AsyncQueue.scala 207:22]
  wire  sourceE_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceE_io_q_sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 207:22]
  wire  sourceE_io_q_sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 207:22]
  wire  sourceE_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 207:22]
  wire  tx_clock; // @[ChipLink.scala 188:20]
  wire  tx_reset; // @[ChipLink.scala 188:20]
  wire  tx_io_c2b_clk; // @[ChipLink.scala 188:20]
  wire  tx_io_c2b_rst; // @[ChipLink.scala 188:20]
  wire  tx_io_c2b_send; // @[ChipLink.scala 188:20]
  wire [7:0] tx_io_c2b_data; // @[ChipLink.scala 188:20]
  wire  tx_io_sa_ready; // @[ChipLink.scala 188:20]
  wire  tx_io_sa_valid; // @[ChipLink.scala 188:20]
  wire [31:0] tx_io_sa_bits_data; // @[ChipLink.scala 188:20]
  wire  tx_io_sa_bits_last; // @[ChipLink.scala 188:20]
  wire [6:0] tx_io_sa_bits_beats; // @[ChipLink.scala 188:20]
  wire  tx_io_sb_ready; // @[ChipLink.scala 188:20]
  wire [31:0] tx_io_sb_bits_data; // @[ChipLink.scala 188:20]
  wire  tx_io_sb_bits_last; // @[ChipLink.scala 188:20]
  wire  tx_io_sc_ready; // @[ChipLink.scala 188:20]
  wire [31:0] tx_io_sc_bits_data; // @[ChipLink.scala 188:20]
  wire  tx_io_sc_bits_last; // @[ChipLink.scala 188:20]
  wire  tx_io_sd_ready; // @[ChipLink.scala 188:20]
  wire  tx_io_sd_valid; // @[ChipLink.scala 188:20]
  wire [31:0] tx_io_sd_bits_data; // @[ChipLink.scala 188:20]
  wire  tx_io_sd_bits_last; // @[ChipLink.scala 188:20]
  wire [6:0] tx_io_sd_bits_beats; // @[ChipLink.scala 188:20]
  wire [31:0] tx_io_se_bits_data; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_rxc_mem_0_a; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_rxc_mem_0_b; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_rxc_mem_0_c; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_rxc_mem_0_d; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_rxc_mem_0_e; // @[ChipLink.scala 188:20]
  wire  tx_io_rxc_ridx; // @[ChipLink.scala 188:20]
  wire  tx_io_rxc_widx; // @[ChipLink.scala 188:20]
  wire  tx_io_rxc_safe_ridx_valid; // @[ChipLink.scala 188:20]
  wire  tx_io_rxc_safe_widx_valid; // @[ChipLink.scala 188:20]
  wire  tx_io_rxc_safe_source_reset_n; // @[ChipLink.scala 188:20]
  wire  tx_io_rxc_safe_sink_reset_n; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_txc_mem_0_a; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_txc_mem_0_b; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_txc_mem_0_c; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_txc_mem_0_d; // @[ChipLink.scala 188:20]
  wire [19:0] tx_io_txc_mem_0_e; // @[ChipLink.scala 188:20]
  wire  tx_io_txc_ridx; // @[ChipLink.scala 188:20]
  wire  tx_io_txc_widx; // @[ChipLink.scala 188:20]
  wire  tx_io_txc_safe_ridx_valid; // @[ChipLink.scala 188:20]
  wire  tx_io_txc_safe_widx_valid; // @[ChipLink.scala 188:20]
  wire  tx_io_txc_safe_source_reset_n; // @[ChipLink.scala 188:20]
  wire  tx_io_txc_safe_sink_reset_n; // @[ChipLink.scala 188:20]
  wire  do_bypass_catcher_clock; // @[ResetCatchAndSync.scala 39:28]
  wire  do_bypass_catcher_reset; // @[ResetCatchAndSync.scala 39:28]
  wire  do_bypass_catcher_io_sync_reset; // @[ResetCatchAndSync.scala 39:28]
  wire  do_bypass_catcher_1_clock; // @[ResetCatchAndSync.scala 39:28]
  wire  do_bypass_catcher_1_reset; // @[ResetCatchAndSync.scala 39:28]
  wire  do_bypass_catcher_1_io_sync_reset; // @[ResetCatchAndSync.scala 39:28]
  TLBusBypass sbypass ( // @[ChipLink.scala 65:35]
    .clock(sbypass_clock),
    .reset(sbypass_reset),
    .auto_node_out_out_a_ready(sbypass_auto_node_out_out_a_ready),
    .auto_node_out_out_a_valid(sbypass_auto_node_out_out_a_valid),
    .auto_node_out_out_a_bits_opcode(sbypass_auto_node_out_out_a_bits_opcode),
    .auto_node_out_out_a_bits_size(sbypass_auto_node_out_out_a_bits_size),
    .auto_node_out_out_a_bits_source(sbypass_auto_node_out_out_a_bits_source),
    .auto_node_out_out_a_bits_address(sbypass_auto_node_out_out_a_bits_address),
    .auto_node_out_out_a_bits_mask(sbypass_auto_node_out_out_a_bits_mask),
    .auto_node_out_out_a_bits_data(sbypass_auto_node_out_out_a_bits_data),
    .auto_node_out_out_d_ready(sbypass_auto_node_out_out_d_ready),
    .auto_node_out_out_d_valid(sbypass_auto_node_out_out_d_valid),
    .auto_node_out_out_d_bits_opcode(sbypass_auto_node_out_out_d_bits_opcode),
    .auto_node_out_out_d_bits_param(sbypass_auto_node_out_out_d_bits_param),
    .auto_node_out_out_d_bits_size(sbypass_auto_node_out_out_d_bits_size),
    .auto_node_out_out_d_bits_source(sbypass_auto_node_out_out_d_bits_source),
    .auto_node_out_out_d_bits_sink(sbypass_auto_node_out_out_d_bits_sink),
    .auto_node_out_out_d_bits_denied(sbypass_auto_node_out_out_d_bits_denied),
    .auto_node_out_out_d_bits_data(sbypass_auto_node_out_out_d_bits_data),
    .auto_node_out_out_d_bits_corrupt(sbypass_auto_node_out_out_d_bits_corrupt),
    .auto_node_in_in_a_ready(sbypass_auto_node_in_in_a_ready),
    .auto_node_in_in_a_valid(sbypass_auto_node_in_in_a_valid),
    .auto_node_in_in_a_bits_opcode(sbypass_auto_node_in_in_a_bits_opcode),
    .auto_node_in_in_a_bits_size(sbypass_auto_node_in_in_a_bits_size),
    .auto_node_in_in_a_bits_source(sbypass_auto_node_in_in_a_bits_source),
    .auto_node_in_in_a_bits_address(sbypass_auto_node_in_in_a_bits_address),
    .auto_node_in_in_a_bits_mask(sbypass_auto_node_in_in_a_bits_mask),
    .auto_node_in_in_a_bits_data(sbypass_auto_node_in_in_a_bits_data),
    .auto_node_in_in_d_ready(sbypass_auto_node_in_in_d_ready),
    .auto_node_in_in_d_valid(sbypass_auto_node_in_in_d_valid),
    .auto_node_in_in_d_bits_opcode(sbypass_auto_node_in_in_d_bits_opcode),
    .auto_node_in_in_d_bits_param(sbypass_auto_node_in_in_d_bits_param),
    .auto_node_in_in_d_bits_size(sbypass_auto_node_in_in_d_bits_size),
    .auto_node_in_in_d_bits_source(sbypass_auto_node_in_in_d_bits_source),
    .auto_node_in_in_d_bits_sink(sbypass_auto_node_in_in_d_bits_sink),
    .auto_node_in_in_d_bits_denied(sbypass_auto_node_in_in_d_bits_denied),
    .auto_node_in_in_d_bits_data(sbypass_auto_node_in_in_d_bits_data),
    .auto_node_in_in_d_bits_corrupt(sbypass_auto_node_in_in_d_bits_corrupt),
    .io_bypass(sbypass_io_bypass)
  );
  StuckSnooper mbypass ( // @[ChipLink.scala 69:35]
    .clock(mbypass_clock),
    .reset(mbypass_reset),
    .auto_in_1_a_ready(mbypass_auto_in_1_a_ready),
    .auto_in_1_a_valid(mbypass_auto_in_1_a_valid),
    .auto_in_1_a_bits_opcode(mbypass_auto_in_1_a_bits_opcode),
    .auto_in_1_a_bits_param(mbypass_auto_in_1_a_bits_param),
    .auto_in_1_a_bits_size(mbypass_auto_in_1_a_bits_size),
    .auto_in_1_a_bits_source(mbypass_auto_in_1_a_bits_source),
    .auto_in_1_a_bits_address(mbypass_auto_in_1_a_bits_address),
    .auto_in_1_a_bits_mask(mbypass_auto_in_1_a_bits_mask),
    .auto_in_1_a_bits_data(mbypass_auto_in_1_a_bits_data),
    .auto_in_1_c_ready(mbypass_auto_in_1_c_ready),
    .auto_in_1_c_valid(mbypass_auto_in_1_c_valid),
    .auto_in_1_c_bits_opcode(mbypass_auto_in_1_c_bits_opcode),
    .auto_in_1_c_bits_param(mbypass_auto_in_1_c_bits_param),
    .auto_in_1_c_bits_size(mbypass_auto_in_1_c_bits_size),
    .auto_in_1_c_bits_source(mbypass_auto_in_1_c_bits_source),
    .auto_in_1_c_bits_address(mbypass_auto_in_1_c_bits_address),
    .auto_in_1_d_ready(mbypass_auto_in_1_d_ready),
    .auto_in_1_d_valid(mbypass_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(mbypass_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_param(mbypass_auto_in_1_d_bits_param),
    .auto_in_1_d_bits_size(mbypass_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_source(mbypass_auto_in_1_d_bits_source),
    .auto_in_1_d_bits_denied(mbypass_auto_in_1_d_bits_denied),
    .auto_in_1_d_bits_data(mbypass_auto_in_1_d_bits_data),
    .auto_in_1_e_ready(mbypass_auto_in_1_e_ready),
    .auto_in_1_e_valid(mbypass_auto_in_1_e_valid),
    .auto_in_1_e_bits_sink(mbypass_auto_in_1_e_bits_sink),
    .auto_out_a_ready(mbypass_auto_out_a_ready),
    .auto_out_a_valid(mbypass_auto_out_a_valid),
    .auto_out_a_bits_opcode(mbypass_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(mbypass_auto_out_a_bits_param),
    .auto_out_a_bits_size(mbypass_auto_out_a_bits_size),
    .auto_out_a_bits_source(mbypass_auto_out_a_bits_source),
    .auto_out_a_bits_address(mbypass_auto_out_a_bits_address),
    .auto_out_a_bits_mask(mbypass_auto_out_a_bits_mask),
    .auto_out_a_bits_data(mbypass_auto_out_a_bits_data),
    .auto_out_c_ready(mbypass_auto_out_c_ready),
    .auto_out_c_valid(mbypass_auto_out_c_valid),
    .auto_out_c_bits_opcode(mbypass_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(mbypass_auto_out_c_bits_param),
    .auto_out_c_bits_size(mbypass_auto_out_c_bits_size),
    .auto_out_c_bits_source(mbypass_auto_out_c_bits_source),
    .auto_out_c_bits_address(mbypass_auto_out_c_bits_address),
    .auto_out_d_ready(mbypass_auto_out_d_ready),
    .auto_out_d_valid(mbypass_auto_out_d_valid),
    .auto_out_d_bits_opcode(mbypass_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(mbypass_auto_out_d_bits_param),
    .auto_out_d_bits_size(mbypass_auto_out_d_bits_size),
    .auto_out_d_bits_source(mbypass_auto_out_d_bits_source),
    .auto_out_d_bits_denied(mbypass_auto_out_d_bits_denied),
    .auto_out_d_bits_data(mbypass_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(mbypass_auto_out_d_bits_corrupt),
    .auto_out_e_ready(mbypass_auto_out_e_ready),
    .auto_out_e_valid(mbypass_auto_out_e_valid),
    .auto_out_e_bits_sink(mbypass_auto_out_e_bits_sink),
    .io_bypass(mbypass_io_bypass)
  );
  TLMonitor_7 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  SinkA sinkA ( // @[ChipLink.scala 148:23]
    .clock(sinkA_clock),
    .reset(sinkA_reset),
    .io_a_ready(sinkA_io_a_ready),
    .io_a_valid(sinkA_io_a_valid),
    .io_a_bits_opcode(sinkA_io_a_bits_opcode),
    .io_a_bits_size(sinkA_io_a_bits_size),
    .io_a_bits_source(sinkA_io_a_bits_source),
    .io_a_bits_address(sinkA_io_a_bits_address),
    .io_a_bits_mask(sinkA_io_a_bits_mask),
    .io_a_bits_data(sinkA_io_a_bits_data),
    .io_q_ready(sinkA_io_q_ready),
    .io_q_valid(sinkA_io_q_valid),
    .io_q_bits_data(sinkA_io_q_bits_data),
    .io_q_bits_last(sinkA_io_q_bits_last),
    .io_q_bits_beats(sinkA_io_q_bits_beats)
  );
  SinkB sinkB ( // @[ChipLink.scala 149:23]
    .clock(sinkB_clock),
    .reset(sinkB_reset),
    .io_q_ready(sinkB_io_q_ready),
    .io_q_valid(sinkB_io_q_valid),
    .io_q_bits_data(sinkB_io_q_bits_data),
    .io_q_bits_last(sinkB_io_q_bits_last)
  );
  SinkC sinkC ( // @[ChipLink.scala 150:23]
    .clock(sinkC_clock),
    .reset(sinkC_reset),
    .io_q_ready(sinkC_io_q_ready),
    .io_q_valid(sinkC_io_q_valid),
    .io_q_bits_data(sinkC_io_q_bits_data),
    .io_q_bits_last(sinkC_io_q_bits_last)
  );
  SinkD sinkD ( // @[ChipLink.scala 151:23]
    .clock(sinkD_clock),
    .reset(sinkD_reset),
    .io_d_ready(sinkD_io_d_ready),
    .io_d_valid(sinkD_io_d_valid),
    .io_d_bits_opcode(sinkD_io_d_bits_opcode),
    .io_d_bits_param(sinkD_io_d_bits_param),
    .io_d_bits_size(sinkD_io_d_bits_size),
    .io_d_bits_source(sinkD_io_d_bits_source),
    .io_d_bits_denied(sinkD_io_d_bits_denied),
    .io_d_bits_data(sinkD_io_d_bits_data),
    .io_q_ready(sinkD_io_q_ready),
    .io_q_valid(sinkD_io_q_valid),
    .io_q_bits_data(sinkD_io_q_bits_data),
    .io_q_bits_last(sinkD_io_q_bits_last),
    .io_q_bits_beats(sinkD_io_q_bits_beats),
    .io_a_tlSource_valid(sinkD_io_a_tlSource_valid),
    .io_a_tlSource_bits(sinkD_io_a_tlSource_bits),
    .io_a_clSource(sinkD_io_a_clSource),
    .io_c_tlSource_valid(sinkD_io_c_tlSource_valid),
    .io_c_tlSource_bits(sinkD_io_c_tlSource_bits),
    .io_c_clSource(sinkD_io_c_clSource)
  );
  SinkE sinkE ( // @[ChipLink.scala 152:23]
    .io_q_bits_data(sinkE_io_q_bits_data),
    .io_d_clSink(sinkE_io_d_clSink)
  );
  SourceA sourceA ( // @[ChipLink.scala 153:25]
    .clock(sourceA_clock),
    .reset(sourceA_reset),
    .io_a_ready(sourceA_io_a_ready),
    .io_a_valid(sourceA_io_a_valid),
    .io_a_bits_opcode(sourceA_io_a_bits_opcode),
    .io_a_bits_param(sourceA_io_a_bits_param),
    .io_a_bits_size(sourceA_io_a_bits_size),
    .io_a_bits_source(sourceA_io_a_bits_source),
    .io_a_bits_address(sourceA_io_a_bits_address),
    .io_a_bits_mask(sourceA_io_a_bits_mask),
    .io_a_bits_data(sourceA_io_a_bits_data),
    .io_q_ready(sourceA_io_q_ready),
    .io_q_valid(sourceA_io_q_valid),
    .io_q_bits(sourceA_io_q_bits),
    .io_d_tlSource_valid(sourceA_io_d_tlSource_valid),
    .io_d_tlSource_bits(sourceA_io_d_tlSource_bits),
    .io_d_clSource(sourceA_io_d_clSource)
  );
  SourceB sourceB ( // @[ChipLink.scala 154:25]
    .clock(sourceB_clock),
    .reset(sourceB_reset),
    .io_q_ready(sourceB_io_q_ready),
    .io_q_valid(sourceB_io_q_valid),
    .io_q_bits(sourceB_io_q_bits)
  );
  SourceC sourceC ( // @[ChipLink.scala 155:25]
    .clock(sourceC_clock),
    .reset(sourceC_reset),
    .io_c_ready(sourceC_io_c_ready),
    .io_c_valid(sourceC_io_c_valid),
    .io_c_bits_opcode(sourceC_io_c_bits_opcode),
    .io_c_bits_param(sourceC_io_c_bits_param),
    .io_c_bits_size(sourceC_io_c_bits_size),
    .io_c_bits_source(sourceC_io_c_bits_source),
    .io_c_bits_address(sourceC_io_c_bits_address),
    .io_q_ready(sourceC_io_q_ready),
    .io_q_valid(sourceC_io_q_valid),
    .io_q_bits(sourceC_io_q_bits),
    .io_d_tlSource_valid(sourceC_io_d_tlSource_valid),
    .io_d_tlSource_bits(sourceC_io_d_tlSource_bits),
    .io_d_clSource(sourceC_io_d_clSource)
  );
  SourceD sourceD ( // @[ChipLink.scala 156:25]
    .clock(sourceD_clock),
    .reset(sourceD_reset),
    .io_d_ready(sourceD_io_d_ready),
    .io_d_valid(sourceD_io_d_valid),
    .io_d_bits_opcode(sourceD_io_d_bits_opcode),
    .io_d_bits_param(sourceD_io_d_bits_param),
    .io_d_bits_size(sourceD_io_d_bits_size),
    .io_d_bits_source(sourceD_io_d_bits_source),
    .io_d_bits_sink(sourceD_io_d_bits_sink),
    .io_d_bits_denied(sourceD_io_d_bits_denied),
    .io_d_bits_data(sourceD_io_d_bits_data),
    .io_d_bits_corrupt(sourceD_io_d_bits_corrupt),
    .io_q_ready(sourceD_io_q_ready),
    .io_q_valid(sourceD_io_q_valid),
    .io_q_bits(sourceD_io_q_bits),
    .io_e_clSink(sourceD_io_e_clSink)
  );
  SourceE sourceE ( // @[ChipLink.scala 157:25]
    .io_e_ready(sourceE_io_e_ready),
    .io_e_valid(sourceE_io_e_valid),
    .io_e_bits_sink(sourceE_io_e_bits_sink),
    .io_q_ready(sourceE_io_q_ready),
    .io_q_valid(sourceE_io_q_valid),
    .io_q_bits(sourceE_io_q_bits)
  );
  RX rx ( // @[ChipLink.scala 159:20]
    .clock(rx_clock),
    .reset(rx_reset),
    .io_b2c_send(rx_io_b2c_send),
    .io_b2c_data(rx_io_b2c_data),
    .io_a_mem_0(rx_io_a_mem_0),
    .io_a_mem_1(rx_io_a_mem_1),
    .io_a_mem_2(rx_io_a_mem_2),
    .io_a_mem_3(rx_io_a_mem_3),
    .io_a_mem_4(rx_io_a_mem_4),
    .io_a_mem_5(rx_io_a_mem_5),
    .io_a_mem_6(rx_io_a_mem_6),
    .io_a_mem_7(rx_io_a_mem_7),
    .io_a_ridx(rx_io_a_ridx),
    .io_a_widx(rx_io_a_widx),
    .io_a_safe_ridx_valid(rx_io_a_safe_ridx_valid),
    .io_a_safe_widx_valid(rx_io_a_safe_widx_valid),
    .io_a_safe_source_reset_n(rx_io_a_safe_source_reset_n),
    .io_a_safe_sink_reset_n(rx_io_a_safe_sink_reset_n),
    .io_bmem_0(rx_io_bmem_0),
    .io_bmem_1(rx_io_bmem_1),
    .io_bmem_2(rx_io_bmem_2),
    .io_bmem_3(rx_io_bmem_3),
    .io_bmem_4(rx_io_bmem_4),
    .io_bmem_5(rx_io_bmem_5),
    .io_bmem_6(rx_io_bmem_6),
    .io_bmem_7(rx_io_bmem_7),
    .io_bridx(rx_io_bridx),
    .io_bwidx(rx_io_bwidx),
    .io_bsafe_ridx_valid(rx_io_bsafe_ridx_valid),
    .io_bsafe_widx_valid(rx_io_bsafe_widx_valid),
    .io_bsafe_source_reset_n(rx_io_bsafe_source_reset_n),
    .io_bsafe_sink_reset_n(rx_io_bsafe_sink_reset_n),
    .io_c_mem_0(rx_io_c_mem_0),
    .io_c_mem_1(rx_io_c_mem_1),
    .io_c_mem_2(rx_io_c_mem_2),
    .io_c_mem_3(rx_io_c_mem_3),
    .io_c_mem_4(rx_io_c_mem_4),
    .io_c_mem_5(rx_io_c_mem_5),
    .io_c_mem_6(rx_io_c_mem_6),
    .io_c_mem_7(rx_io_c_mem_7),
    .io_c_ridx(rx_io_c_ridx),
    .io_c_widx(rx_io_c_widx),
    .io_c_safe_ridx_valid(rx_io_c_safe_ridx_valid),
    .io_c_safe_widx_valid(rx_io_c_safe_widx_valid),
    .io_c_safe_source_reset_n(rx_io_c_safe_source_reset_n),
    .io_c_safe_sink_reset_n(rx_io_c_safe_sink_reset_n),
    .io_d_mem_0(rx_io_d_mem_0),
    .io_d_mem_1(rx_io_d_mem_1),
    .io_d_mem_2(rx_io_d_mem_2),
    .io_d_mem_3(rx_io_d_mem_3),
    .io_d_mem_4(rx_io_d_mem_4),
    .io_d_mem_5(rx_io_d_mem_5),
    .io_d_mem_6(rx_io_d_mem_6),
    .io_d_mem_7(rx_io_d_mem_7),
    .io_d_ridx(rx_io_d_ridx),
    .io_d_widx(rx_io_d_widx),
    .io_d_safe_ridx_valid(rx_io_d_safe_ridx_valid),
    .io_d_safe_widx_valid(rx_io_d_safe_widx_valid),
    .io_d_safe_source_reset_n(rx_io_d_safe_source_reset_n),
    .io_d_safe_sink_reset_n(rx_io_d_safe_sink_reset_n),
    .io_e_mem_0(rx_io_e_mem_0),
    .io_e_mem_1(rx_io_e_mem_1),
    .io_e_mem_2(rx_io_e_mem_2),
    .io_e_mem_3(rx_io_e_mem_3),
    .io_e_mem_4(rx_io_e_mem_4),
    .io_e_mem_5(rx_io_e_mem_5),
    .io_e_mem_6(rx_io_e_mem_6),
    .io_e_mem_7(rx_io_e_mem_7),
    .io_e_ridx(rx_io_e_ridx),
    .io_e_widx(rx_io_e_widx),
    .io_e_safe_ridx_valid(rx_io_e_safe_ridx_valid),
    .io_e_safe_widx_valid(rx_io_e_safe_widx_valid),
    .io_e_safe_source_reset_n(rx_io_e_safe_source_reset_n),
    .io_e_safe_sink_reset_n(rx_io_e_safe_sink_reset_n),
    .io_rxc_mem_0_a(rx_io_rxc_mem_0_a),
    .io_rxc_mem_0_b(rx_io_rxc_mem_0_b),
    .io_rxc_mem_0_c(rx_io_rxc_mem_0_c),
    .io_rxc_mem_0_d(rx_io_rxc_mem_0_d),
    .io_rxc_mem_0_e(rx_io_rxc_mem_0_e),
    .io_rxc_ridx(rx_io_rxc_ridx),
    .io_rxc_widx(rx_io_rxc_widx),
    .io_rxc_safe_ridx_valid(rx_io_rxc_safe_ridx_valid),
    .io_rxc_safe_widx_valid(rx_io_rxc_safe_widx_valid),
    .io_rxc_safe_source_reset_n(rx_io_rxc_safe_source_reset_n),
    .io_rxc_safe_sink_reset_n(rx_io_rxc_safe_sink_reset_n),
    .io_txc_mem_0_a(rx_io_txc_mem_0_a),
    .io_txc_mem_0_b(rx_io_txc_mem_0_b),
    .io_txc_mem_0_c(rx_io_txc_mem_0_c),
    .io_txc_mem_0_d(rx_io_txc_mem_0_d),
    .io_txc_mem_0_e(rx_io_txc_mem_0_e),
    .io_txc_ridx(rx_io_txc_ridx),
    .io_txc_widx(rx_io_txc_widx),
    .io_txc_safe_ridx_valid(rx_io_txc_safe_ridx_valid),
    .io_txc_safe_widx_valid(rx_io_txc_safe_widx_valid),
    .io_txc_safe_source_reset_n(rx_io_txc_safe_source_reset_n),
    .io_txc_safe_sink_reset_n(rx_io_txc_safe_sink_reset_n)
  );
  AsyncResetReg rx_reset_reg ( // @[AsyncResetReg.scala 74:21]
    .io_q(rx_reset_reg_io_q),
    .io_clk(rx_reset_reg_io_clk),
    .io_rst(rx_reset_reg_io_rst)
  );
  AsyncQueueSink sourceA_io_q_sink ( // @[AsyncQueue.scala 207:22]
    .clock(sourceA_io_q_sink_clock),
    .reset(sourceA_io_q_sink_reset),
    .io_deq_ready(sourceA_io_q_sink_io_deq_ready),
    .io_deq_valid(sourceA_io_q_sink_io_deq_valid),
    .io_deq_bits(sourceA_io_q_sink_io_deq_bits),
    .io_async_mem_0(sourceA_io_q_sink_io_async_mem_0),
    .io_async_mem_1(sourceA_io_q_sink_io_async_mem_1),
    .io_async_mem_2(sourceA_io_q_sink_io_async_mem_2),
    .io_async_mem_3(sourceA_io_q_sink_io_async_mem_3),
    .io_async_mem_4(sourceA_io_q_sink_io_async_mem_4),
    .io_async_mem_5(sourceA_io_q_sink_io_async_mem_5),
    .io_async_mem_6(sourceA_io_q_sink_io_async_mem_6),
    .io_async_mem_7(sourceA_io_q_sink_io_async_mem_7),
    .io_async_ridx(sourceA_io_q_sink_io_async_ridx),
    .io_async_widx(sourceA_io_q_sink_io_async_widx),
    .io_async_safe_ridx_valid(sourceA_io_q_sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(sourceA_io_q_sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(sourceA_io_q_sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(sourceA_io_q_sink_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink sourceB_io_q_sink ( // @[AsyncQueue.scala 207:22]
    .clock(sourceB_io_q_sink_clock),
    .reset(sourceB_io_q_sink_reset),
    .io_deq_ready(sourceB_io_q_sink_io_deq_ready),
    .io_deq_valid(sourceB_io_q_sink_io_deq_valid),
    .io_deq_bits(sourceB_io_q_sink_io_deq_bits),
    .io_async_mem_0(sourceB_io_q_sink_io_async_mem_0),
    .io_async_mem_1(sourceB_io_q_sink_io_async_mem_1),
    .io_async_mem_2(sourceB_io_q_sink_io_async_mem_2),
    .io_async_mem_3(sourceB_io_q_sink_io_async_mem_3),
    .io_async_mem_4(sourceB_io_q_sink_io_async_mem_4),
    .io_async_mem_5(sourceB_io_q_sink_io_async_mem_5),
    .io_async_mem_6(sourceB_io_q_sink_io_async_mem_6),
    .io_async_mem_7(sourceB_io_q_sink_io_async_mem_7),
    .io_async_ridx(sourceB_io_q_sink_io_async_ridx),
    .io_async_widx(sourceB_io_q_sink_io_async_widx),
    .io_async_safe_ridx_valid(sourceB_io_q_sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(sourceB_io_q_sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(sourceB_io_q_sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(sourceB_io_q_sink_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink sourceC_io_q_sink ( // @[AsyncQueue.scala 207:22]
    .clock(sourceC_io_q_sink_clock),
    .reset(sourceC_io_q_sink_reset),
    .io_deq_ready(sourceC_io_q_sink_io_deq_ready),
    .io_deq_valid(sourceC_io_q_sink_io_deq_valid),
    .io_deq_bits(sourceC_io_q_sink_io_deq_bits),
    .io_async_mem_0(sourceC_io_q_sink_io_async_mem_0),
    .io_async_mem_1(sourceC_io_q_sink_io_async_mem_1),
    .io_async_mem_2(sourceC_io_q_sink_io_async_mem_2),
    .io_async_mem_3(sourceC_io_q_sink_io_async_mem_3),
    .io_async_mem_4(sourceC_io_q_sink_io_async_mem_4),
    .io_async_mem_5(sourceC_io_q_sink_io_async_mem_5),
    .io_async_mem_6(sourceC_io_q_sink_io_async_mem_6),
    .io_async_mem_7(sourceC_io_q_sink_io_async_mem_7),
    .io_async_ridx(sourceC_io_q_sink_io_async_ridx),
    .io_async_widx(sourceC_io_q_sink_io_async_widx),
    .io_async_safe_ridx_valid(sourceC_io_q_sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(sourceC_io_q_sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(sourceC_io_q_sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(sourceC_io_q_sink_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink sourceD_io_q_sink ( // @[AsyncQueue.scala 207:22]
    .clock(sourceD_io_q_sink_clock),
    .reset(sourceD_io_q_sink_reset),
    .io_deq_ready(sourceD_io_q_sink_io_deq_ready),
    .io_deq_valid(sourceD_io_q_sink_io_deq_valid),
    .io_deq_bits(sourceD_io_q_sink_io_deq_bits),
    .io_async_mem_0(sourceD_io_q_sink_io_async_mem_0),
    .io_async_mem_1(sourceD_io_q_sink_io_async_mem_1),
    .io_async_mem_2(sourceD_io_q_sink_io_async_mem_2),
    .io_async_mem_3(sourceD_io_q_sink_io_async_mem_3),
    .io_async_mem_4(sourceD_io_q_sink_io_async_mem_4),
    .io_async_mem_5(sourceD_io_q_sink_io_async_mem_5),
    .io_async_mem_6(sourceD_io_q_sink_io_async_mem_6),
    .io_async_mem_7(sourceD_io_q_sink_io_async_mem_7),
    .io_async_ridx(sourceD_io_q_sink_io_async_ridx),
    .io_async_widx(sourceD_io_q_sink_io_async_widx),
    .io_async_safe_ridx_valid(sourceD_io_q_sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(sourceD_io_q_sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(sourceD_io_q_sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(sourceD_io_q_sink_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink sourceE_io_q_sink ( // @[AsyncQueue.scala 207:22]
    .clock(sourceE_io_q_sink_clock),
    .reset(sourceE_io_q_sink_reset),
    .io_deq_ready(sourceE_io_q_sink_io_deq_ready),
    .io_deq_valid(sourceE_io_q_sink_io_deq_valid),
    .io_deq_bits(sourceE_io_q_sink_io_deq_bits),
    .io_async_mem_0(sourceE_io_q_sink_io_async_mem_0),
    .io_async_mem_1(sourceE_io_q_sink_io_async_mem_1),
    .io_async_mem_2(sourceE_io_q_sink_io_async_mem_2),
    .io_async_mem_3(sourceE_io_q_sink_io_async_mem_3),
    .io_async_mem_4(sourceE_io_q_sink_io_async_mem_4),
    .io_async_mem_5(sourceE_io_q_sink_io_async_mem_5),
    .io_async_mem_6(sourceE_io_q_sink_io_async_mem_6),
    .io_async_mem_7(sourceE_io_q_sink_io_async_mem_7),
    .io_async_ridx(sourceE_io_q_sink_io_async_ridx),
    .io_async_widx(sourceE_io_q_sink_io_async_widx),
    .io_async_safe_ridx_valid(sourceE_io_q_sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(sourceE_io_q_sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(sourceE_io_q_sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(sourceE_io_q_sink_io_async_safe_sink_reset_n)
  );
  TX tx ( // @[ChipLink.scala 188:20]
    .clock(tx_clock),
    .reset(tx_reset),
    .io_c2b_clk(tx_io_c2b_clk),
    .io_c2b_rst(tx_io_c2b_rst),
    .io_c2b_send(tx_io_c2b_send),
    .io_c2b_data(tx_io_c2b_data),
    .io_sa_ready(tx_io_sa_ready),
    .io_sa_valid(tx_io_sa_valid),
    .io_sa_bits_data(tx_io_sa_bits_data),
    .io_sa_bits_last(tx_io_sa_bits_last),
    .io_sa_bits_beats(tx_io_sa_bits_beats),
    .io_sb_ready(tx_io_sb_ready),
    .io_sb_bits_data(tx_io_sb_bits_data),
    .io_sb_bits_last(tx_io_sb_bits_last),
    .io_sc_ready(tx_io_sc_ready),
    .io_sc_bits_data(tx_io_sc_bits_data),
    .io_sc_bits_last(tx_io_sc_bits_last),
    .io_sd_ready(tx_io_sd_ready),
    .io_sd_valid(tx_io_sd_valid),
    .io_sd_bits_data(tx_io_sd_bits_data),
    .io_sd_bits_last(tx_io_sd_bits_last),
    .io_sd_bits_beats(tx_io_sd_bits_beats),
    .io_se_bits_data(tx_io_se_bits_data),
    .io_rxc_mem_0_a(tx_io_rxc_mem_0_a),
    .io_rxc_mem_0_b(tx_io_rxc_mem_0_b),
    .io_rxc_mem_0_c(tx_io_rxc_mem_0_c),
    .io_rxc_mem_0_d(tx_io_rxc_mem_0_d),
    .io_rxc_mem_0_e(tx_io_rxc_mem_0_e),
    .io_rxc_ridx(tx_io_rxc_ridx),
    .io_rxc_widx(tx_io_rxc_widx),
    .io_rxc_safe_ridx_valid(tx_io_rxc_safe_ridx_valid),
    .io_rxc_safe_widx_valid(tx_io_rxc_safe_widx_valid),
    .io_rxc_safe_source_reset_n(tx_io_rxc_safe_source_reset_n),
    .io_rxc_safe_sink_reset_n(tx_io_rxc_safe_sink_reset_n),
    .io_txc_mem_0_a(tx_io_txc_mem_0_a),
    .io_txc_mem_0_b(tx_io_txc_mem_0_b),
    .io_txc_mem_0_c(tx_io_txc_mem_0_c),
    .io_txc_mem_0_d(tx_io_txc_mem_0_d),
    .io_txc_mem_0_e(tx_io_txc_mem_0_e),
    .io_txc_ridx(tx_io_txc_ridx),
    .io_txc_widx(tx_io_txc_widx),
    .io_txc_safe_ridx_valid(tx_io_txc_safe_ridx_valid),
    .io_txc_safe_widx_valid(tx_io_txc_safe_widx_valid),
    .io_txc_safe_source_reset_n(tx_io_txc_safe_source_reset_n),
    .io_txc_safe_sink_reset_n(tx_io_txc_safe_sink_reset_n)
  );
  ResetCatchAndSync_d3 do_bypass_catcher ( // @[ResetCatchAndSync.scala 39:28]
    .clock(do_bypass_catcher_clock),
    .reset(do_bypass_catcher_reset),
    .io_sync_reset(do_bypass_catcher_io_sync_reset)
  );
  ResetCatchAndSync_d3 do_bypass_catcher_1 ( // @[ResetCatchAndSync.scala 39:28]
    .clock(do_bypass_catcher_1_clock),
    .reset(do_bypass_catcher_1_reset),
    .io_sync_reset(do_bypass_catcher_1_io_sync_reset)
  );
  assign auto_mbypass_out_a_valid = mbypass_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_a_bits_opcode = mbypass_auto_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_a_bits_param = mbypass_auto_out_a_bits_param; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_a_bits_size = mbypass_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_a_bits_source = mbypass_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_a_bits_address = mbypass_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_a_bits_mask = mbypass_auto_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_a_bits_data = mbypass_auto_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_c_valid = mbypass_auto_out_c_valid; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_c_bits_opcode = mbypass_auto_out_c_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_c_bits_param = mbypass_auto_out_c_bits_param; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_c_bits_size = mbypass_auto_out_c_bits_size; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_c_bits_source = mbypass_auto_out_c_bits_source; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_c_bits_address = mbypass_auto_out_c_bits_address; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_d_ready = mbypass_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_e_valid = mbypass_auto_out_e_valid; // @[LazyModule.scala 311:12]
  assign auto_mbypass_out_e_bits_sink = mbypass_auto_out_e_bits_sink; // @[LazyModule.scala 311:12]
  assign auto_sbypass_node_in_in_a_ready = sbypass_auto_node_in_in_a_ready; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_valid = sbypass_auto_node_in_in_d_valid; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_bits_opcode = sbypass_auto_node_in_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_bits_param = sbypass_auto_node_in_in_d_bits_param; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_bits_size = sbypass_auto_node_in_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_bits_source = sbypass_auto_node_in_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_bits_sink = sbypass_auto_node_in_in_d_bits_sink; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_bits_denied = sbypass_auto_node_in_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_bits_data = sbypass_auto_node_in_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign auto_sbypass_node_in_in_d_bits_corrupt = sbypass_auto_node_in_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign auto_io_out_c2b_clk = tx_io_c2b_clk; // @[Nodes.scala 1207:84 ChipLink.scala 189:18]
  assign auto_io_out_c2b_rst = tx_io_c2b_rst; // @[Nodes.scala 1207:84 ChipLink.scala 190:18]
  assign auto_io_out_c2b_send = tx_io_c2b_send; // @[Nodes.scala 1207:84 ChipLink.scala 192:19]
  assign auto_io_out_c2b_data = tx_io_c2b_data; // @[Nodes.scala 1207:84 ChipLink.scala 191:19]
  assign sbypass_clock = clock;
  assign sbypass_reset = reset;
  assign sbypass_auto_node_out_out_a_ready = sinkA_io_a_ready; // @[Nodes.scala 1210:84 ChipLink.scala 193:16]
  assign sbypass_auto_node_out_out_d_valid = sourceD_io_d_valid; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_out_out_d_bits_opcode = sourceD_io_d_bits_opcode; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_out_out_d_bits_param = sourceD_io_d_bits_param; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_out_out_d_bits_size = sourceD_io_d_bits_size; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_out_out_d_bits_source = sourceD_io_d_bits_source; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_out_out_d_bits_sink = sourceD_io_d_bits_sink; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_out_out_d_bits_denied = sourceD_io_d_bits_denied; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_out_out_d_bits_data = sourceD_io_d_bits_data; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_out_out_d_bits_corrupt = sourceD_io_d_bits_corrupt; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sbypass_auto_node_in_in_a_valid = auto_sbypass_node_in_in_a_valid; // @[LazyModule.scala 309:16]
  assign sbypass_auto_node_in_in_a_bits_opcode = auto_sbypass_node_in_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign sbypass_auto_node_in_in_a_bits_size = auto_sbypass_node_in_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign sbypass_auto_node_in_in_a_bits_source = auto_sbypass_node_in_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign sbypass_auto_node_in_in_a_bits_address = auto_sbypass_node_in_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign sbypass_auto_node_in_in_a_bits_mask = auto_sbypass_node_in_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign sbypass_auto_node_in_in_a_bits_data = auto_sbypass_node_in_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign sbypass_auto_node_in_in_d_ready = auto_sbypass_node_in_in_d_ready; // @[LazyModule.scala 309:16]
  assign sbypass_io_bypass = do_bypass_catcher_io_sync_reset | do_bypass_catcher_1_io_sync_reset; // @[ChipLink.scala 228:56]
  assign mbypass_clock = clock;
  assign mbypass_reset = reset;
  assign mbypass_auto_in_1_a_valid = sourceA_io_a_valid; // @[Nodes.scala 1207:84 ChipLink.scala 177:11]
  assign mbypass_auto_in_1_a_bits_opcode = sourceA_io_a_bits_opcode; // @[Nodes.scala 1207:84 ChipLink.scala 177:11]
  assign mbypass_auto_in_1_a_bits_param = sourceA_io_a_bits_param; // @[Nodes.scala 1207:84 ChipLink.scala 177:11]
  assign mbypass_auto_in_1_a_bits_size = sourceA_io_a_bits_size; // @[Nodes.scala 1207:84 ChipLink.scala 177:11]
  assign mbypass_auto_in_1_a_bits_source = sourceA_io_a_bits_source; // @[Nodes.scala 1207:84 ChipLink.scala 177:11]
  assign mbypass_auto_in_1_a_bits_address = sourceA_io_a_bits_address; // @[Nodes.scala 1207:84 ChipLink.scala 177:11]
  assign mbypass_auto_in_1_a_bits_mask = sourceA_io_a_bits_mask; // @[Nodes.scala 1207:84 ChipLink.scala 177:11]
  assign mbypass_auto_in_1_a_bits_data = sourceA_io_a_bits_data; // @[Nodes.scala 1207:84 ChipLink.scala 177:11]
  assign mbypass_auto_in_1_c_valid = sourceC_io_c_valid; // @[Nodes.scala 1207:84 ChipLink.scala 179:11]
  assign mbypass_auto_in_1_c_bits_opcode = sourceC_io_c_bits_opcode; // @[Nodes.scala 1207:84 ChipLink.scala 179:11]
  assign mbypass_auto_in_1_c_bits_param = sourceC_io_c_bits_param; // @[Nodes.scala 1207:84 ChipLink.scala 179:11]
  assign mbypass_auto_in_1_c_bits_size = sourceC_io_c_bits_size; // @[Nodes.scala 1207:84 ChipLink.scala 179:11]
  assign mbypass_auto_in_1_c_bits_source = sourceC_io_c_bits_source; // @[Nodes.scala 1207:84 ChipLink.scala 179:11]
  assign mbypass_auto_in_1_c_bits_address = sourceC_io_c_bits_address; // @[Nodes.scala 1207:84 ChipLink.scala 179:11]
  assign mbypass_auto_in_1_d_ready = sinkD_io_d_ready; // @[Nodes.scala 1207:84 ChipLink.scala 196:16]
  assign mbypass_auto_in_1_e_valid = sourceE_io_e_valid; // @[Nodes.scala 1207:84 ChipLink.scala 181:11]
  assign mbypass_auto_in_1_e_bits_sink = sourceE_io_e_bits_sink; // @[Nodes.scala 1207:84 ChipLink.scala 181:11]
  assign mbypass_auto_out_a_ready = auto_mbypass_out_a_ready; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_c_ready = auto_mbypass_out_c_ready; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_d_valid = auto_mbypass_out_d_valid; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_d_bits_opcode = auto_mbypass_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_d_bits_param = auto_mbypass_out_d_bits_param; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_d_bits_size = auto_mbypass_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_d_bits_source = auto_mbypass_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_d_bits_denied = auto_mbypass_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_d_bits_data = auto_mbypass_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_d_bits_corrupt = auto_mbypass_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign mbypass_auto_out_e_ready = auto_mbypass_out_e_ready; // @[LazyModule.scala 311:12]
  assign mbypass_io_bypass = do_bypass_catcher_io_sync_reset | do_bypass_catcher_1_io_sync_reset; // @[ChipLink.scala 228:56]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = sinkA_io_a_ready; // @[Nodes.scala 1210:84 ChipLink.scala 193:16]
  assign monitor_io_in_a_valid = sbypass_auto_node_out_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign monitor_io_in_a_bits_opcode = sbypass_auto_node_out_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign monitor_io_in_a_bits_size = sbypass_auto_node_out_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign monitor_io_in_a_bits_source = sbypass_auto_node_out_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign monitor_io_in_a_bits_address = sbypass_auto_node_out_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign monitor_io_in_a_bits_mask = sbypass_auto_node_out_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign monitor_io_in_d_ready = sbypass_auto_node_out_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign monitor_io_in_d_valid = sourceD_io_d_valid; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign monitor_io_in_d_bits_opcode = sourceD_io_d_bits_opcode; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign monitor_io_in_d_bits_param = sourceD_io_d_bits_param; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign monitor_io_in_d_bits_size = sourceD_io_d_bits_size; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign monitor_io_in_d_bits_source = sourceD_io_d_bits_source; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign monitor_io_in_d_bits_sink = sourceD_io_d_bits_sink; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign monitor_io_in_d_bits_denied = sourceD_io_d_bits_denied; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign monitor_io_in_d_bits_corrupt = sourceD_io_d_bits_corrupt; // @[Nodes.scala 1210:84 ChipLink.scala 180:11]
  assign sinkA_clock = clock;
  assign sinkA_reset = reset;
  assign sinkA_io_a_valid = sbypass_auto_node_out_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign sinkA_io_a_bits_opcode = sbypass_auto_node_out_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign sinkA_io_a_bits_size = sbypass_auto_node_out_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign sinkA_io_a_bits_source = sbypass_auto_node_out_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign sinkA_io_a_bits_address = sbypass_auto_node_out_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign sinkA_io_a_bits_mask = sbypass_auto_node_out_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign sinkA_io_a_bits_data = sbypass_auto_node_out_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign sinkA_io_q_ready = tx_io_sa_ready; // @[ChipLink.scala 199:16]
  assign sinkB_clock = clock;
  assign sinkB_reset = reset;
  assign sinkB_io_q_ready = tx_io_sb_ready; // @[ChipLink.scala 200:16]
  assign sinkC_clock = clock;
  assign sinkC_reset = reset;
  assign sinkC_io_q_ready = tx_io_sc_ready; // @[ChipLink.scala 201:16]
  assign sinkD_clock = clock;
  assign sinkD_reset = reset;
  assign sinkD_io_d_valid = mbypass_auto_in_1_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sinkD_io_d_bits_opcode = mbypass_auto_in_1_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sinkD_io_d_bits_param = mbypass_auto_in_1_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sinkD_io_d_bits_size = mbypass_auto_in_1_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sinkD_io_d_bits_source = mbypass_auto_in_1_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sinkD_io_d_bits_denied = mbypass_auto_in_1_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sinkD_io_d_bits_data = mbypass_auto_in_1_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sinkD_io_q_ready = tx_io_sd_ready; // @[ChipLink.scala 202:16]
  assign sinkD_io_a_clSource = sourceA_io_d_clSource; // @[ChipLink.scala 220:25]
  assign sinkD_io_c_clSource = sourceC_io_d_clSource; // @[ChipLink.scala 222:25]
  assign sinkE_io_d_clSink = sourceD_io_e_clSink; // @[ChipLink.scala 225:23]
  assign sourceA_clock = clock;
  assign sourceA_reset = reset;
  assign sourceA_io_a_ready = mbypass_auto_in_1_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sourceA_io_q_valid = sourceA_io_q_sink_io_deq_valid; // @[ChipLink.scala 182:18]
  assign sourceA_io_q_bits = sourceA_io_q_sink_io_deq_bits; // @[ChipLink.scala 182:18]
  assign sourceA_io_d_tlSource_valid = sinkD_io_a_tlSource_valid; // @[ChipLink.scala 221:27]
  assign sourceA_io_d_tlSource_bits = sinkD_io_a_tlSource_bits; // @[ChipLink.scala 221:27]
  assign sourceB_clock = clock;
  assign sourceB_reset = reset;
  assign sourceB_io_q_valid = sourceB_io_q_sink_io_deq_valid; // @[ChipLink.scala 183:18]
  assign sourceB_io_q_bits = sourceB_io_q_sink_io_deq_bits; // @[ChipLink.scala 183:18]
  assign sourceC_clock = clock;
  assign sourceC_reset = reset;
  assign sourceC_io_c_ready = mbypass_auto_in_1_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sourceC_io_q_valid = sourceC_io_q_sink_io_deq_valid; // @[ChipLink.scala 184:18]
  assign sourceC_io_q_bits = sourceC_io_q_sink_io_deq_bits; // @[ChipLink.scala 184:18]
  assign sourceC_io_d_tlSource_valid = sinkD_io_c_tlSource_valid; // @[ChipLink.scala 223:27]
  assign sourceC_io_d_tlSource_bits = sinkD_io_c_tlSource_bits; // @[ChipLink.scala 223:27]
  assign sourceD_clock = clock;
  assign sourceD_reset = reset;
  assign sourceD_io_d_ready = sbypass_auto_node_out_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign sourceD_io_q_valid = sourceD_io_q_sink_io_deq_valid; // @[ChipLink.scala 185:18]
  assign sourceD_io_q_bits = sourceD_io_q_sink_io_deq_bits; // @[ChipLink.scala 185:18]
  assign sourceE_io_e_ready = mbypass_auto_in_1_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign sourceE_io_q_valid = sourceE_io_q_sink_io_deq_valid; // @[ChipLink.scala 186:18]
  assign sourceE_io_q_bits = sourceE_io_q_sink_io_deq_bits; // @[ChipLink.scala 186:18]
  assign rx_clock = auto_io_out_b2c_clk; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign rx_reset = rx_reset_reg_io_q; // @[ChipLink.scala 168:18]
  assign rx_io_b2c_send = auto_io_out_b2c_send; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign rx_io_b2c_data = auto_io_out_b2c_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign rx_io_a_ridx = sourceA_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 208:19]
  assign rx_io_a_safe_ridx_valid = sourceA_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 208:19]
  assign rx_io_a_safe_sink_reset_n = sourceA_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 208:19]
  assign rx_io_bridx = sourceB_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 208:19]
  assign rx_io_bsafe_ridx_valid = sourceB_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 208:19]
  assign rx_io_bsafe_sink_reset_n = sourceB_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 208:19]
  assign rx_io_c_ridx = sourceC_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 208:19]
  assign rx_io_c_safe_ridx_valid = sourceC_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 208:19]
  assign rx_io_c_safe_sink_reset_n = sourceC_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 208:19]
  assign rx_io_d_ridx = sourceD_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 208:19]
  assign rx_io_d_safe_ridx_valid = sourceD_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 208:19]
  assign rx_io_d_safe_sink_reset_n = sourceD_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 208:19]
  assign rx_io_e_ridx = sourceE_io_q_sink_io_async_ridx; // @[AsyncQueue.scala 208:19]
  assign rx_io_e_safe_ridx_valid = sourceE_io_q_sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 208:19]
  assign rx_io_e_safe_sink_reset_n = sourceE_io_q_sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 208:19]
  assign rx_io_rxc_ridx = tx_io_rxc_ridx; // @[ChipLink.scala 216:15]
  assign rx_io_rxc_safe_ridx_valid = tx_io_rxc_safe_ridx_valid; // @[ChipLink.scala 216:15]
  assign rx_io_rxc_safe_sink_reset_n = tx_io_rxc_safe_sink_reset_n; // @[ChipLink.scala 216:15]
  assign rx_io_txc_ridx = tx_io_txc_ridx; // @[ChipLink.scala 217:15]
  assign rx_io_txc_safe_ridx_valid = tx_io_txc_safe_ridx_valid; // @[ChipLink.scala 217:15]
  assign rx_io_txc_safe_sink_reset_n = tx_io_txc_safe_sink_reset_n; // @[ChipLink.scala 217:15]
  assign rx_reset_reg_io_clk = auto_io_out_b2c_clk; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign rx_reset_reg_io_rst = auto_io_out_b2c_rst; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign sourceA_io_q_sink_clock = clock;
  assign sourceA_io_q_sink_reset = reset;
  assign sourceA_io_q_sink_io_deq_ready = sourceA_io_q_ready; // @[ChipLink.scala 182:18]
  assign sourceA_io_q_sink_io_async_mem_0 = rx_io_a_mem_0; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_mem_1 = rx_io_a_mem_1; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_mem_2 = rx_io_a_mem_2; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_mem_3 = rx_io_a_mem_3; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_mem_4 = rx_io_a_mem_4; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_mem_5 = rx_io_a_mem_5; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_mem_6 = rx_io_a_mem_6; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_mem_7 = rx_io_a_mem_7; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_widx = rx_io_a_widx; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_safe_widx_valid = rx_io_a_safe_widx_valid; // @[AsyncQueue.scala 208:19]
  assign sourceA_io_q_sink_io_async_safe_source_reset_n = rx_io_a_safe_source_reset_n; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_clock = clock;
  assign sourceB_io_q_sink_reset = reset;
  assign sourceB_io_q_sink_io_deq_ready = sourceB_io_q_ready; // @[ChipLink.scala 183:18]
  assign sourceB_io_q_sink_io_async_mem_0 = rx_io_bmem_0; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_mem_1 = rx_io_bmem_1; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_mem_2 = rx_io_bmem_2; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_mem_3 = rx_io_bmem_3; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_mem_4 = rx_io_bmem_4; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_mem_5 = rx_io_bmem_5; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_mem_6 = rx_io_bmem_6; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_mem_7 = rx_io_bmem_7; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_widx = rx_io_bwidx; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_safe_widx_valid = rx_io_bsafe_widx_valid; // @[AsyncQueue.scala 208:19]
  assign sourceB_io_q_sink_io_async_safe_source_reset_n = rx_io_bsafe_source_reset_n; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_clock = clock;
  assign sourceC_io_q_sink_reset = reset;
  assign sourceC_io_q_sink_io_deq_ready = sourceC_io_q_ready; // @[ChipLink.scala 184:18]
  assign sourceC_io_q_sink_io_async_mem_0 = rx_io_c_mem_0; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_mem_1 = rx_io_c_mem_1; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_mem_2 = rx_io_c_mem_2; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_mem_3 = rx_io_c_mem_3; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_mem_4 = rx_io_c_mem_4; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_mem_5 = rx_io_c_mem_5; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_mem_6 = rx_io_c_mem_6; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_mem_7 = rx_io_c_mem_7; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_widx = rx_io_c_widx; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_safe_widx_valid = rx_io_c_safe_widx_valid; // @[AsyncQueue.scala 208:19]
  assign sourceC_io_q_sink_io_async_safe_source_reset_n = rx_io_c_safe_source_reset_n; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_clock = clock;
  assign sourceD_io_q_sink_reset = reset;
  assign sourceD_io_q_sink_io_deq_ready = sourceD_io_q_ready; // @[ChipLink.scala 185:18]
  assign sourceD_io_q_sink_io_async_mem_0 = rx_io_d_mem_0; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_mem_1 = rx_io_d_mem_1; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_mem_2 = rx_io_d_mem_2; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_mem_3 = rx_io_d_mem_3; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_mem_4 = rx_io_d_mem_4; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_mem_5 = rx_io_d_mem_5; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_mem_6 = rx_io_d_mem_6; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_mem_7 = rx_io_d_mem_7; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_widx = rx_io_d_widx; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_safe_widx_valid = rx_io_d_safe_widx_valid; // @[AsyncQueue.scala 208:19]
  assign sourceD_io_q_sink_io_async_safe_source_reset_n = rx_io_d_safe_source_reset_n; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_clock = clock;
  assign sourceE_io_q_sink_reset = reset;
  assign sourceE_io_q_sink_io_deq_ready = sourceE_io_q_ready; // @[ChipLink.scala 186:18]
  assign sourceE_io_q_sink_io_async_mem_0 = rx_io_e_mem_0; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_mem_1 = rx_io_e_mem_1; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_mem_2 = rx_io_e_mem_2; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_mem_3 = rx_io_e_mem_3; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_mem_4 = rx_io_e_mem_4; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_mem_5 = rx_io_e_mem_5; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_mem_6 = rx_io_e_mem_6; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_mem_7 = rx_io_e_mem_7; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_widx = rx_io_e_widx; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_safe_widx_valid = rx_io_e_safe_widx_valid; // @[AsyncQueue.scala 208:19]
  assign sourceE_io_q_sink_io_async_safe_source_reset_n = rx_io_e_safe_source_reset_n; // @[AsyncQueue.scala 208:19]
  assign tx_clock = clock;
  assign tx_reset = reset;
  assign tx_io_sa_valid = sinkA_io_q_valid; // @[ChipLink.scala 199:16]
  assign tx_io_sa_bits_data = sinkA_io_q_bits_data; // @[ChipLink.scala 199:16]
  assign tx_io_sa_bits_last = sinkA_io_q_bits_last; // @[ChipLink.scala 199:16]
  assign tx_io_sa_bits_beats = sinkA_io_q_bits_beats; // @[ChipLink.scala 199:16]
  assign tx_io_sb_bits_data = sinkB_io_q_bits_data; // @[ChipLink.scala 200:16]
  assign tx_io_sb_bits_last = sinkB_io_q_bits_last; // @[ChipLink.scala 200:16]
  assign tx_io_sc_bits_data = sinkC_io_q_bits_data; // @[ChipLink.scala 201:16]
  assign tx_io_sc_bits_last = sinkC_io_q_bits_last; // @[ChipLink.scala 201:16]
  assign tx_io_sd_valid = sinkD_io_q_valid; // @[ChipLink.scala 202:16]
  assign tx_io_sd_bits_data = sinkD_io_q_bits_data; // @[ChipLink.scala 202:16]
  assign tx_io_sd_bits_last = sinkD_io_q_bits_last; // @[ChipLink.scala 202:16]
  assign tx_io_sd_bits_beats = sinkD_io_q_bits_beats; // @[ChipLink.scala 202:16]
  assign tx_io_se_bits_data = sinkE_io_q_bits_data; // @[ChipLink.scala 203:16]
  assign tx_io_rxc_mem_0_a = rx_io_rxc_mem_0_a; // @[ChipLink.scala 216:15]
  assign tx_io_rxc_mem_0_b = rx_io_rxc_mem_0_b; // @[ChipLink.scala 216:15]
  assign tx_io_rxc_mem_0_c = rx_io_rxc_mem_0_c; // @[ChipLink.scala 216:15]
  assign tx_io_rxc_mem_0_d = rx_io_rxc_mem_0_d; // @[ChipLink.scala 216:15]
  assign tx_io_rxc_mem_0_e = rx_io_rxc_mem_0_e; // @[ChipLink.scala 216:15]
  assign tx_io_rxc_widx = rx_io_rxc_widx; // @[ChipLink.scala 216:15]
  assign tx_io_rxc_safe_widx_valid = rx_io_rxc_safe_widx_valid; // @[ChipLink.scala 216:15]
  assign tx_io_rxc_safe_source_reset_n = rx_io_rxc_safe_source_reset_n; // @[ChipLink.scala 216:15]
  assign tx_io_txc_mem_0_a = rx_io_txc_mem_0_a; // @[ChipLink.scala 217:15]
  assign tx_io_txc_mem_0_b = rx_io_txc_mem_0_b; // @[ChipLink.scala 217:15]
  assign tx_io_txc_mem_0_c = rx_io_txc_mem_0_c; // @[ChipLink.scala 217:15]
  assign tx_io_txc_mem_0_d = rx_io_txc_mem_0_d; // @[ChipLink.scala 217:15]
  assign tx_io_txc_mem_0_e = rx_io_txc_mem_0_e; // @[ChipLink.scala 217:15]
  assign tx_io_txc_widx = rx_io_txc_widx; // @[ChipLink.scala 217:15]
  assign tx_io_txc_safe_widx_valid = rx_io_txc_safe_widx_valid; // @[ChipLink.scala 217:15]
  assign tx_io_txc_safe_source_reset_n = rx_io_txc_safe_source_reset_n; // @[ChipLink.scala 217:15]
  assign do_bypass_catcher_clock = clock;
  assign do_bypass_catcher_reset = rx_reset; // @[compatibility.scala 260:56]
  assign do_bypass_catcher_1_clock = clock;
  assign do_bypass_catcher_1_reset = tx_reset; // @[compatibility.scala 260:56]
endmodule
module TLMonitor_8(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [3:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [3:0]  io_in_a_bits_mask,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [3:0]  io_in_d_bits_source,
  input  [5:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = ~io_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | io_in_a_bits_source[3]; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_34 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_60 = 3'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48]
  wire [31:0] _T_62 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_63 = {1'b0,$signed(_T_62)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_65 = $signed(_T_63) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_66 = $signed(_T_65) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_77 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_78 = {1'b0,$signed(_T_77)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_80 = $signed(_T_78) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_81 = $signed(_T_80) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_82 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_83 = {1'b0,$signed(_T_82)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_85 = $signed(_T_83) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_86 = $signed(_T_85) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_90 = _T_66 | _T_71 | _T_76 | _T_81 | _T_86; // @[Parameters.scala 671:42]
  wire  _T_91 = _T_60 & _T_90; // @[Parameters.scala 670:56]
  wire  _T_93 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_96 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_97 = {1'b0,$signed(_T_96)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_99 = $signed(_T_97) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_100 = $signed(_T_99) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_101 = _T_93 & _T_100; // @[Parameters.scala 670:56]
  wire  _T_104 = _T_91 | _T_101; // @[Parameters.scala 672:30]
  wire  _T_105 = source_ok & _T_104; // @[Monitor.scala 82:72]
  wire [32:0] _T_136 = $signed(_T_78) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _T_137 = $signed(_T_136) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_141 = _T_100 | _T_66 | _T_71 | _T_76 | _T_137; // @[Parameters.scala 671:42]
  wire [3:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_163 = _T_162 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_312 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_367 = _T_93 & _T_141; // @[Parameters.scala 670:56]
  wire  _T_382 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_390 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_444 = source_ok & _T_367; // @[Monitor.scala 115:71]
  wire  _T_462 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_530 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_531 = io_in_a_bits_mask & _T_530; // @[Monitor.scala 127:31]
  wire  _T_532 = _T_531 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_536 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_556 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_581 = _T_66 | _T_71 | _T_76 | _T_137; // @[Parameters.scala 671:42]
  wire  _T_582 = _T_556 & _T_581; // @[Parameters.scala 670:56]
  wire  _T_594 = _T_582 | _T_101; // @[Parameters.scala 672:30]
  wire  _T_595 = source_ok & _T_594; // @[Monitor.scala 131:74]
  wire  _T_613 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_690 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_766 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_13 = ~io_in_d_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_13 | io_in_d_bits_source[3]; // @[Parameters.scala 1125:46]
  wire  sink_ok = io_in_d_bits_sink < 6'h21; // @[Monitor.scala 306:31]
  wire  _T_770 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_774 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_778 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_782 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_786 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_790 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_801 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_805 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_818 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_838 = _T_786 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_847 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_864 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_882 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [3:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_912 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_913 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_921 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_925 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_929 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [3:0] source_1; // @[Monitor.scala 538:22]
  reg [5:0] sink; // @[Monitor.scala 539:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_936 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_937 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_941 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_945 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_949 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_953 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29]
  wire  _T_957 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [15:0] inflight; // @[Monitor.scala 611:27]
  reg [63:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [63:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69]
  wire [63:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [63:0] _GEN_73 = {{48'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[63:1]}; // @[Monitor.scala 634:152]
  wire [63:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [63:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91]
  wire [63:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[63:1]}; // @[Monitor.scala 638:144]
  wire  _T_963 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire  _T_966 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [15:0] _T_968 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_970 = ~_T_968[0]; // @[Monitor.scala 658:17]
  wire [15:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [130:0] _GEN_19 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [130:0] _GEN_20 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_974 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_976 = ~_T_770; // @[Monitor.scala 671:74]
  wire  _T_977 = io_in_d_valid & d_first_1 & ~_T_770; // @[Monitor.scala 671:71]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [15:0] d_clr = _d_first_T & d_first_1 & _T_976 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [142:0] _GEN_23 = _d_first_T & d_first_1 & _T_976 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_963 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [15:0] _T_987 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_989 = _T_987[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_994 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39]
  wire  _T_995 = io_in_d_bits_opcode == _GEN_32 | _T_994; // @[Monitor.scala 685:77]
  wire  _T_999 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_1006 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_1007 = io_in_d_bits_opcode == _GEN_48 | _T_1006; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_1011 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_1021 = _T_974 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_976; // @[Monitor.scala 694:116]
  wire  _T_1023 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire [15:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [15:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [15:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [63:0] a_opcodes_set = _GEN_19[63:0];
  wire [63:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [63:0] d_opcodes_clr = _GEN_23[63:0];
  wire [63:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [63:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [63:0] a_sizes_set = _GEN_20[63:0];
  wire [63:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [63:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_1032 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [15:0] inflight_1; // @[Monitor.scala 723:35]
  reg [63:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [63:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [63:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93]
  wire [63:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[63:1]}; // @[Monitor.scala 747:146]
  wire  _T_1058 = io_in_d_valid & d_first_2 & _T_770; // @[Monitor.scala 779:71]
  wire [15:0] d_clr_1 = _d_first_T & d_first_2 & _T_770 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [142:0] _GEN_68 = _d_first_T & d_first_2 & _T_770 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire [15:0] _T_1066 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_1076 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [15:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [15:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [63:0] d_opcodes_clr_1 = _GEN_68[63:0];
  wire [63:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [63:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_1096 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 16'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 64'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 64'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 16'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 64'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_105 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_105 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_163 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_163 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_105 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_105 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_163 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_163 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_367 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_367 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_532 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_532 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_595 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_595 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_595 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_595 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_766 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_766 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_786 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_786 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(sink_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(sink_ok | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_801 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_805 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(sink_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(sink_ok | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_801 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_805 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_838 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_838 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_838 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_838 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_913 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_913 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_921 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_921 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_925 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_925 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_929 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_929 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_937 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_937 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_941 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_941 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_945 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_945 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_949 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_949 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_953 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_953 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_957 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_957 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_966 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_966 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~(_T_989 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~(_T_989 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_995 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_995 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_999 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_999 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1007 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1007 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1011 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1011 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1021 & ~(_T_1023 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1021 & ~(_T_1023 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1032 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1032 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1058 & ~(_T_1066[0] | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1058 & ~(_T_1066[0] | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1058 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1058 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1096 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:102:43)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1096 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  source = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  address = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  d_first_counter = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  opcode_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  param_1 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  sink = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight = _RAND_12[15:0];
  _RAND_13 = {2{`RANDOM}};
  inflight_opcodes = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_sizes = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  watchdog = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  inflight_1 = _RAND_18[15:0];
  _RAND_19 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  watchdog_1 = _RAND_21[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFIFOFixer(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [3:0]  auto_in_a_bits_mask,
  input  [31:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output [5:0]  auto_in_d_bits_sink,
  output        auto_in_d_bits_denied,
  output [31:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [3:0]  auto_out_a_bits_mask,
  output [31:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [2:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input  [5:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [31:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire [32:0] _a_notFIFO_T_1 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T = auto_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_1 = {1'b0,$signed(_a_id_T)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_3 = $signed(_a_id_T_1) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_4 = $signed(_a_id_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _a_id_T_5 = auto_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_6 = {1'b0,$signed(_a_id_T_5)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_8 = $signed(_a_id_T_6) & 33'she0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_9 = $signed(_a_id_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _a_id_T_10 = auto_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_11 = {1'b0,$signed(_a_id_T_10)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_13 = $signed(_a_id_T_11) & 33'shc0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_14 = $signed(_a_id_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _a_id_T_15 = auto_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_16 = {1'b0,$signed(_a_id_T_15)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_18 = $signed(_a_id_T_16) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_19 = $signed(_a_id_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _a_id_T_22 = _a_id_T_4 | _a_id_T_9 | _a_id_T_14 | _a_id_T_19; // @[Parameters.scala 615:89]
  wire [32:0] _a_id_T_26 = $signed(_a_notFIFO_T_1) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_27 = $signed(_a_id_T_26) == 33'sh0; // @[Parameters.scala 137:67]
  wire [1:0] _a_id_T_29 = _a_id_T_27 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_70 = {{1'd0}, _a_id_T_22}; // @[Mux.scala 27:72]
  wire [1:0] a_id = _GEN_70 | _a_id_T_29; // @[Mux.scala 27:72]
  wire  a_noDomain = a_id == 2'h0; // @[FIFOFixer.scala 55:29]
  wire  stalls_a_sel = ~auto_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg  flight_0; // @[FIFOFixer.scala 71:27]
  reg  flight_1; // @[FIFOFixer.scala 71:27]
  reg  flight_2; // @[FIFOFixer.scala 71:27]
  reg  flight_3; // @[FIFOFixer.scala 71:27]
  reg  flight_4; // @[FIFOFixer.scala 71:27]
  reg  flight_5; // @[FIFOFixer.scala 71:27]
  reg  flight_6; // @[FIFOFixer.scala 71:27]
  reg  flight_7; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id; // @[Reg.scala 15:16]
  wire  stalls_0 = stalls_a_sel & a_first & (flight_0 | flight_1 | flight_2 | flight_3 | flight_4 | flight_5 | flight_6
     | flight_7) & (a_noDomain | stalls_id != a_id); // @[FIFOFixer.scala 80:50]
  reg  flight_8; // @[FIFOFixer.scala 71:27]
  reg  flight_9; // @[FIFOFixer.scala 71:27]
  reg  flight_10; // @[FIFOFixer.scala 71:27]
  reg  flight_11; // @[FIFOFixer.scala 71:27]
  reg  flight_12; // @[FIFOFixer.scala 71:27]
  reg  flight_13; // @[FIFOFixer.scala 71:27]
  reg  flight_14; // @[FIFOFixer.scala 71:27]
  reg  flight_15; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id_1; // @[Reg.scala 15:16]
  wire  stalls_1 = auto_in_a_bits_source[3] & a_first & (flight_8 | flight_9 | flight_10 | flight_11 | flight_12 |
    flight_13 | flight_14 | flight_15) & (a_noDomain | stalls_id_1 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stall = stalls_0 | stalls_1; // @[FIFOFixer.scala 83:49]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[FIFOFixer.scala 88:50]
  wire  bundleIn_0_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  wire  _a_first_T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _a_first_beats1_decode_T_1 = 13'h3f << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _a_first_beats1_decode_T_3 = ~_a_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] a_first_beats1_decode = _a_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  _d_first_T = auto_in_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  wire  d_first = d_first_first & auto_out_d_bits_opcode != 3'h6; // @[FIFOFixer.scala 67:42]
  wire  _GEN_18 = a_first & _a_first_T ? 4'h0 == auto_in_a_bits_source | flight_0 : flight_0; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_19 = a_first & _a_first_T ? 4'h1 == auto_in_a_bits_source | flight_1 : flight_1; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_20 = a_first & _a_first_T ? 4'h2 == auto_in_a_bits_source | flight_2 : flight_2; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_21 = a_first & _a_first_T ? 4'h3 == auto_in_a_bits_source | flight_3 : flight_3; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_22 = a_first & _a_first_T ? 4'h4 == auto_in_a_bits_source | flight_4 : flight_4; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_23 = a_first & _a_first_T ? 4'h5 == auto_in_a_bits_source | flight_5 : flight_5; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_24 = a_first & _a_first_T ? 4'h6 == auto_in_a_bits_source | flight_6 : flight_6; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_25 = a_first & _a_first_T ? 4'h7 == auto_in_a_bits_source | flight_7 : flight_7; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_26 = a_first & _a_first_T ? 4'h8 == auto_in_a_bits_source | flight_8 : flight_8; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_27 = a_first & _a_first_T ? 4'h9 == auto_in_a_bits_source | flight_9 : flight_9; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_28 = a_first & _a_first_T ? 4'ha == auto_in_a_bits_source | flight_10 : flight_10; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_29 = a_first & _a_first_T ? 4'hb == auto_in_a_bits_source | flight_11 : flight_11; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_30 = a_first & _a_first_T ? 4'hc == auto_in_a_bits_source | flight_12 : flight_12; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_31 = a_first & _a_first_T ? 4'hd == auto_in_a_bits_source | flight_13 : flight_13; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_32 = a_first & _a_first_T ? 4'he == auto_in_a_bits_source | flight_14 : flight_14; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_33 = a_first & _a_first_T ? 4'hf == auto_in_a_bits_source | flight_15 : flight_15; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _stalls_id_T_1 = _a_first_T & stalls_a_sel; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_5 = _a_first_T & auto_in_a_bits_source[3]; // @[FIFOFixer.scala 77:49]
  TLMonitor_8 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  assign auto_in_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  assign auto_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid & _bundleIn_0_a_ready_T; // @[FIFOFixer.scala 87:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_0 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h0 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_0 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_0 <= _GEN_18;
      end
    end else begin
      flight_0 <= _GEN_18;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_1 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h1 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_1 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_1 <= _GEN_19;
      end
    end else begin
      flight_1 <= _GEN_19;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_2 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h2 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_2 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_2 <= _GEN_20;
      end
    end else begin
      flight_2 <= _GEN_20;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_3 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h3 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_3 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_3 <= _GEN_21;
      end
    end else begin
      flight_3 <= _GEN_21;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_4 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h4 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_4 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_4 <= _GEN_22;
      end
    end else begin
      flight_4 <= _GEN_22;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_5 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h5 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_5 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_5 <= _GEN_23;
      end
    end else begin
      flight_5 <= _GEN_23;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_6 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h6 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_6 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_6 <= _GEN_24;
      end
    end else begin
      flight_6 <= _GEN_24;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_7 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h7 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_7 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_7 <= _GEN_25;
      end
    end else begin
      flight_7 <= _GEN_25;
    end
    if (_stalls_id_T_1) begin // @[Reg.scala 16:19]
      stalls_id <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_8 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h8 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_8 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_8 <= _GEN_26;
      end
    end else begin
      flight_8 <= _GEN_26;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_9 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'h9 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_9 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_9 <= _GEN_27;
      end
    end else begin
      flight_9 <= _GEN_27;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_10 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'ha == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_10 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_10 <= _GEN_28;
      end
    end else begin
      flight_10 <= _GEN_28;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_11 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'hb == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_11 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_11 <= _GEN_29;
      end
    end else begin
      flight_11 <= _GEN_29;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_12 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'hc == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_12 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_12 <= _GEN_30;
      end
    end else begin
      flight_12 <= _GEN_30;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_13 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'hd == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_13 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_13 <= _GEN_31;
      end
    end else begin
      flight_13 <= _GEN_31;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_14 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'he == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_14 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_14 <= _GEN_32;
      end
    end else begin
      flight_14 <= _GEN_32;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_15 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (4'hf == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_15 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_15 <= _GEN_33;
      end
    end else begin
      flight_15 <= _GEN_33;
    end
    if (_stalls_id_T_5) begin // @[Reg.scala 16:19]
      stalls_id_1 <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  flight_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  flight_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  flight_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  flight_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  flight_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  flight_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  flight_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  flight_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  stalls_id = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  flight_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  flight_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  flight_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  flight_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  flight_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  flight_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  flight_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  flight_15 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  stalls_id_1 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  d_first_counter = _RAND_19[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_9(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [3:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [3:0]  io_in_d_bits_source,
  input  [5:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = ~io_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | io_in_a_bits_source[3]; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_2 = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_3 = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_4 = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_5 = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_lo = mask_acc_2 | mask_size_2 & mask_eq_6; // @[Misc.scala 214:29]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_hi = mask_acc_2 | mask_size_2 & mask_eq_7; // @[Misc.scala 214:29]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_lo = mask_acc_3 | mask_size_2 & mask_eq_8; // @[Misc.scala 214:29]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_hi = mask_acc_3 | mask_size_2 & mask_eq_9; // @[Misc.scala 214:29]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_lo = mask_acc_4 | mask_size_2 & mask_eq_10; // @[Misc.scala 214:29]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_hi = mask_acc_4 | mask_size_2 & mask_eq_11; // @[Misc.scala 214:29]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_lo = mask_acc_5 | mask_size_2 & mask_eq_12; // @[Misc.scala 214:29]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_hi = mask_acc_5 | mask_size_2 & mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_34 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_60 = 3'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48]
  wire [31:0] _T_62 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_63 = {1'b0,$signed(_T_62)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_65 = $signed(_T_63) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_66 = $signed(_T_65) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_77 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_78 = {1'b0,$signed(_T_77)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_80 = $signed(_T_78) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_81 = $signed(_T_80) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_82 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_83 = {1'b0,$signed(_T_82)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_85 = $signed(_T_83) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_86 = $signed(_T_85) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_90 = _T_66 | _T_71 | _T_76 | _T_81 | _T_86; // @[Parameters.scala 671:42]
  wire  _T_91 = _T_60 & _T_90; // @[Parameters.scala 670:56]
  wire  _T_93 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_96 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_97 = {1'b0,$signed(_T_96)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_99 = $signed(_T_97) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_100 = $signed(_T_99) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_101 = _T_93 & _T_100; // @[Parameters.scala 670:56]
  wire  _T_104 = _T_91 | _T_101; // @[Parameters.scala 672:30]
  wire  _T_105 = source_ok & _T_104; // @[Monitor.scala 82:72]
  wire [32:0] _T_136 = $signed(_T_78) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _T_137 = $signed(_T_136) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_141 = _T_100 | _T_66 | _T_71 | _T_76 | _T_137; // @[Parameters.scala 671:42]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_312 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_367 = _T_93 & _T_141; // @[Parameters.scala 670:56]
  wire  _T_382 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_390 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_444 = source_ok & _T_367; // @[Monitor.scala 115:71]
  wire  _T_462 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [7:0] _T_530 = ~mask; // @[Monitor.scala 127:33]
  wire [7:0] _T_531 = io_in_a_bits_mask & _T_530; // @[Monitor.scala 127:31]
  wire  _T_532 = _T_531 == 8'h0; // @[Monitor.scala 127:40]
  wire  _T_536 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_556 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_581 = _T_66 | _T_71 | _T_76 | _T_137; // @[Parameters.scala 671:42]
  wire  _T_582 = _T_556 & _T_581; // @[Parameters.scala 670:56]
  wire  _T_594 = _T_582 | _T_101; // @[Parameters.scala 672:30]
  wire  _T_595 = source_ok & _T_594; // @[Monitor.scala 131:74]
  wire  _T_613 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_690 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_766 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_13 = ~io_in_d_bits_source[3]; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_13 | io_in_d_bits_source[3]; // @[Parameters.scala 1125:46]
  wire  sink_ok = io_in_d_bits_sink < 6'h21; // @[Monitor.scala 306:31]
  wire  _T_770 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_774 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27]
  wire  _T_778 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_782 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_786 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_790 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_801 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_805 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_818 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_838 = _T_786 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_847 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_864 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_882 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [3:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_912 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_913 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_921 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_925 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_929 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [3:0] source_1; // @[Monitor.scala 538:22]
  reg [5:0] sink; // @[Monitor.scala 539:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_936 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_937 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_941 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_945 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_949 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_953 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29]
  wire  _T_957 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [15:0] inflight; // @[Monitor.scala 611:27]
  reg [63:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [63:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69]
  wire [63:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [63:0] _GEN_73 = {{48'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97]
  wire [63:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[63:1]}; // @[Monitor.scala 634:152]
  wire [63:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [63:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91]
  wire [63:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[63:1]}; // @[Monitor.scala 638:144]
  wire  _T_963 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire  _T_966 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [15:0] _T_968 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_970 = ~_T_968[0]; // @[Monitor.scala 658:17]
  wire [15:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [130:0] _GEN_19 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [130:0] _GEN_20 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_974 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_976 = ~_T_770; // @[Monitor.scala 671:74]
  wire  _T_977 = io_in_d_valid & d_first_1 & ~_T_770; // @[Monitor.scala 671:71]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [15:0] d_clr = _d_first_T & d_first_1 & _T_976 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [142:0] _GEN_23 = _d_first_T & d_first_1 & _T_976 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_963 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [15:0] _T_987 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_989 = _T_987[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_994 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39]
  wire  _T_995 = io_in_d_bits_opcode == _GEN_32 | _T_994; // @[Monitor.scala 685:77]
  wire  _T_999 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_1006 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_1007 = io_in_d_bits_opcode == _GEN_48 | _T_1006; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_1011 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_1021 = _T_974 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_976; // @[Monitor.scala 694:116]
  wire  _T_1023 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire [15:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [15:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [15:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [63:0] a_opcodes_set = _GEN_19[63:0];
  wire [63:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [63:0] d_opcodes_clr = _GEN_23[63:0];
  wire [63:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [63:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [63:0] a_sizes_set = _GEN_20[63:0];
  wire [63:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [63:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_1032 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [15:0] inflight_1; // @[Monitor.scala 723:35]
  reg [63:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25]
  wire [63:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [63:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93]
  wire [63:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[63:1]}; // @[Monitor.scala 747:146]
  wire  _T_1058 = io_in_d_valid & d_first_2 & _T_770; // @[Monitor.scala 779:71]
  wire [15:0] d_clr_1 = _d_first_T & d_first_2 & _T_770 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [142:0] _GEN_68 = _d_first_T & d_first_2 & _T_770 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire [15:0] _T_1066 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_1076 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [15:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [15:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [63:0] d_opcodes_clr_1 = _GEN_68[63:0];
  wire [63:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [63:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_1096 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 16'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 64'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 64'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 16'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 64'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_105 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_105 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_163 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_34 & ~(_T_163 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_105 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_105 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_163 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & ~(_T_163 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_367 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_367 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_312 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_532 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_462 & ~(_T_532 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_595 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_595 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_536 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_595 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_595 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_613 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_444 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_444 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_382 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_690 & ~(_T_382 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_766 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_766 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_786 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_770 & ~(_T_786 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(sink_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(sink_ok | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_801 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_805 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_790 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(sink_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(sink_ok | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_774 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_774 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_801 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_805 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_838 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_818 & ~(_T_838 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_847 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_838 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_864 & ~(_T_838 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_778 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_778 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_782 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_882 & ~(_T_782 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_913 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_913 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_921 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_921 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_925 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_925 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~(_T_929 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~(_T_929 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_937 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_937 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_941 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_941 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_945 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_945 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_949 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_949 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_953 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_953 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~(_T_957 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~(_T_957 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_966 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_966 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~(_T_989 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~(_T_989 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_995 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_995 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_999 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & same_cycle_resp & ~(_T_999 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1007 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1007 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1011 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~same_cycle_resp & ~(_T_1011 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1021 & ~(_T_1023 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1021 & ~(_T_1023 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1032 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1032 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1058 & ~(_T_1066[0] | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1058 & ~(_T_1066[0] | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1058 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1058 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1096 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:103:7)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1096 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  source = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  address = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  d_first_counter = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  opcode_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  param_1 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  sink = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight = _RAND_12[15:0];
  _RAND_13 = {2{`RANDOM}};
  inflight_opcodes = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_sizes = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  watchdog = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  inflight_1 = _RAND_18[15:0];
  _RAND_19 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  watchdog_1 = _RAND_21[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [3:0] saved_source; // @[Repeater.scala 20:18]
  reg [31:0] saved_address; // @[Repeater.scala 20:18]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18]
  reg [63:0] saved_data; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 28:38 Repeater.scala 28:45 Repeater.scala 19:21]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign io_deq_bits_data = full ? saved_data : io_enq_bits_data; // @[Repeater.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin // @[Repeater.scala 29:38]
      full <= 1'h0; // @[Repeater.scala 29:45]
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_data <= io_enq_bits_data; // @[Repeater.scala 28:62]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_source = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  saved_address = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  saved_mask = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  saved_data = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLWidthWidget(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [3:0]  auto_out_a_bits_mask,
  output [31:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [2:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input  [5:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [31:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  repeated_repeater_clock; // @[Repeater.scala 35:26]
  wire  repeated_repeater_reset; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_repeat; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_size; // @[Repeater.scala 35:26]
  wire [3:0] repeated_repeater_io_enq_bits_source; // @[Repeater.scala 35:26]
  wire [31:0] repeated_repeater_io_enq_bits_address; // @[Repeater.scala 35:26]
  wire [7:0] repeated_repeater_io_enq_bits_mask; // @[Repeater.scala 35:26]
  wire [63:0] repeated_repeater_io_enq_bits_data; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_size; // @[Repeater.scala 35:26]
  wire [3:0] repeated_repeater_io_deq_bits_source; // @[Repeater.scala 35:26]
  wire [31:0] repeated_repeater_io_deq_bits_address; // @[Repeater.scala 35:26]
  wire [7:0] repeated_repeater_io_deq_bits_mask; // @[Repeater.scala 35:26]
  wire [63:0] repeated_repeater_io_deq_bits_data; // @[Repeater.scala 35:26]
  wire [31:0] cated_bits_data_hi = repeated_repeater_io_deq_bits_data[63:32]; // @[WidthWidget.scala 158:37]
  wire [31:0] cated_bits_data_lo = auto_in_a_bits_data[31:0]; // @[WidthWidget.scala 159:31]
  wire [63:0] cated_bits_data = {cated_bits_data_hi,cated_bits_data_lo}; // @[Cat.scala 30:58]
  wire [2:0] cated_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  repeat_hasData = ~cated_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] cated_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire [9:0] _repeat_limit_T_1 = 10'h7 << cated_bits_size; // @[package.scala 234:77]
  wire [2:0] _repeat_limit_T_3 = ~_repeat_limit_T_1[2:0]; // @[package.scala 234:46]
  wire  repeat_limit = _repeat_limit_T_3[2]; // @[WidthWidget.scala 97:47]
  reg  repeat_count; // @[WidthWidget.scala 99:26]
  wire  repeat_last = repeat_count == repeat_limit | ~repeat_hasData; // @[WidthWidget.scala 101:35]
  wire  cated_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  _repeat_T = auto_out_a_ready & cated_valid; // @[Decoupled.scala 40:37]
  wire [31:0] cated_bits_address = repeated_repeater_io_deq_bits_address; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  repeat_sel = cated_bits_address[2]; // @[WidthWidget.scala 110:39]
  wire  repeat_index = repeat_sel | repeat_count; // @[WidthWidget.scala 120:24]
  wire [31:0] repeat_bundleOut_0_a_bits_data_mux_0 = cated_bits_data[31:0]; // @[WidthWidget.scala 122:55]
  wire [31:0] repeat_bundleOut_0_a_bits_data_mux_1 = cated_bits_data[63:32]; // @[WidthWidget.scala 122:55]
  wire [7:0] cated_bits_mask = repeated_repeater_io_deq_bits_mask; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire [3:0] repeat_bundleOut_0_a_bits_mask_mux_0 = cated_bits_mask[3:0]; // @[WidthWidget.scala 122:55]
  wire [3:0] repeat_bundleOut_0_a_bits_mask_mux_1 = cated_bits_mask[7:4]; // @[WidthWidget.scala 122:55]
  wire  hasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [9:0] _limit_T_1 = 10'h7 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [2:0] _limit_T_3 = ~_limit_T_1[2:0]; // @[package.scala 234:46]
  wire  limit = _limit_T_3[2]; // @[WidthWidget.scala 32:47]
  reg  count; // @[WidthWidget.scala 34:27]
  wire  last = count == limit | ~hasData; // @[WidthWidget.scala 36:36]
  wire  enable_0 = ~(|(count & limit)); // @[WidthWidget.scala 37:47]
  reg  corrupt_reg; // @[WidthWidget.scala 39:32]
  wire  corrupt_out = auto_out_d_bits_corrupt | corrupt_reg; // @[WidthWidget.scala 41:36]
  wire  _bundleOut_0_d_ready_T = ~last; // @[WidthWidget.scala 70:32]
  wire  bundleOut_0_d_ready = auto_in_d_ready | ~last; // @[WidthWidget.scala 70:29]
  wire  _T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  reg  bundleIn_0_d_bits_data_rdata_written_once; // @[WidthWidget.scala 56:41]
  wire  bundleIn_0_d_bits_data_masked_enable_0 = enable_0 | ~bundleIn_0_d_bits_data_rdata_written_once; // @[WidthWidget.scala 57:42]
  reg [31:0] bundleIn_0_d_bits_data_rdata_0; // @[WidthWidget.scala 60:24]
  wire [31:0] bundleIn_0_d_bits_data_lo = bundleIn_0_d_bits_data_masked_enable_0 ? auto_out_d_bits_data :
    bundleIn_0_d_bits_data_rdata_0; // @[WidthWidget.scala 62:88]
  wire  _GEN_10 = _T & _bundleOut_0_d_ready_T | bundleIn_0_d_bits_data_rdata_written_once; // @[WidthWidget.scala 63:35 WidthWidget.scala 64:30 WidthWidget.scala 56:41]
  TLMonitor_9 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Repeater repeated_repeater ( // @[Repeater.scala 35:26]
    .clock(repeated_repeater_clock),
    .reset(repeated_repeater_reset),
    .io_repeat(repeated_repeater_io_repeat),
    .io_enq_ready(repeated_repeater_io_enq_ready),
    .io_enq_valid(repeated_repeater_io_enq_valid),
    .io_enq_bits_opcode(repeated_repeater_io_enq_bits_opcode),
    .io_enq_bits_size(repeated_repeater_io_enq_bits_size),
    .io_enq_bits_source(repeated_repeater_io_enq_bits_source),
    .io_enq_bits_address(repeated_repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeated_repeater_io_enq_bits_mask),
    .io_enq_bits_data(repeated_repeater_io_enq_bits_data),
    .io_deq_ready(repeated_repeater_io_deq_ready),
    .io_deq_valid(repeated_repeater_io_deq_valid),
    .io_deq_bits_opcode(repeated_repeater_io_deq_bits_opcode),
    .io_deq_bits_size(repeated_repeater_io_deq_bits_size),
    .io_deq_bits_source(repeated_repeater_io_deq_bits_source),
    .io_deq_bits_address(repeated_repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeated_repeater_io_deq_bits_mask),
    .io_deq_bits_data(repeated_repeater_io_deq_bits_data)
  );
  assign auto_in_a_ready = repeated_repeater_io_enq_ready; // @[Nodes.scala 1210:84 Repeater.scala 37:21]
  assign auto_in_d_valid = auto_out_d_valid & last; // @[WidthWidget.scala 71:29]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = {auto_out_d_bits_data,bundleIn_0_d_bits_data_lo}; // @[Cat.scala 30:58]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt | corrupt_reg; // @[WidthWidget.scala 41:36]
  assign auto_out_a_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_source = repeated_repeater_io_deq_bits_source; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_address = repeated_repeater_io_deq_bits_address; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_mask = repeat_index ? repeat_bundleOut_0_a_bits_mask_mux_1 :
    repeat_bundleOut_0_a_bits_mask_mux_0; // @[WidthWidget.scala 134:53 WidthWidget.scala 134:53]
  assign auto_out_a_bits_data = repeat_index ? repeat_bundleOut_0_a_bits_data_mux_1 :
    repeat_bundleOut_0_a_bits_data_mux_0; // @[WidthWidget.scala 131:30 WidthWidget.scala 131:30]
  assign auto_out_d_ready = auto_in_d_ready | ~last; // @[WidthWidget.scala 70:29]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = repeated_repeater_io_enq_ready; // @[Nodes.scala 1210:84 Repeater.scala 37:21]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = auto_out_d_valid & last; // @[WidthWidget.scala 71:29]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt | corrupt_reg; // @[WidthWidget.scala 41:36]
  assign repeated_repeater_clock = clock;
  assign repeated_repeater_reset = reset;
  assign repeated_repeater_io_repeat = ~repeat_last; // @[WidthWidget.scala 142:7]
  assign repeated_repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  always @(posedge clock) begin
    if (reset) begin // @[WidthWidget.scala 99:26]
      repeat_count <= 1'h0; // @[WidthWidget.scala 99:26]
    end else if (_repeat_T) begin // @[WidthWidget.scala 103:25]
      if (repeat_last) begin // @[WidthWidget.scala 105:21]
        repeat_count <= 1'h0; // @[WidthWidget.scala 105:29]
      end else begin
        repeat_count <= repeat_count + 1'h1; // @[WidthWidget.scala 104:15]
      end
    end
    if (reset) begin // @[WidthWidget.scala 34:27]
      count <= 1'h0; // @[WidthWidget.scala 34:27]
    end else if (_T) begin // @[WidthWidget.scala 43:24]
      if (last) begin // @[WidthWidget.scala 46:21]
        count <= 1'h0; // @[WidthWidget.scala 47:17]
      end else begin
        count <= count + 1'h1; // @[WidthWidget.scala 44:15]
      end
    end
    if (reset) begin // @[WidthWidget.scala 39:32]
      corrupt_reg <= 1'h0; // @[WidthWidget.scala 39:32]
    end else if (_T) begin // @[WidthWidget.scala 43:24]
      if (last) begin // @[WidthWidget.scala 46:21]
        corrupt_reg <= 1'h0; // @[WidthWidget.scala 48:23]
      end else begin
        corrupt_reg <= corrupt_out; // @[WidthWidget.scala 45:21]
      end
    end
    if (reset) begin // @[WidthWidget.scala 56:41]
      bundleIn_0_d_bits_data_rdata_written_once <= 1'h0; // @[WidthWidget.scala 56:41]
    end else begin
      bundleIn_0_d_bits_data_rdata_written_once <= _GEN_10;
    end
    if (_T & _bundleOut_0_d_ready_T) begin // @[WidthWidget.scala 63:35]
      if (bundleIn_0_d_bits_data_masked_enable_0) begin // @[WidthWidget.scala 62:88]
        bundleIn_0_d_bits_data_rdata_0 <= auto_out_d_bits_data;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  repeat_count = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  corrupt_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bundleIn_0_d_bits_data_rdata_written_once = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bundleIn_0_d_bits_data_rdata_0 = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_11(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ram_id [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_resp [0:0]; // @[Decoupled.scala 218:16]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_last [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_10 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 249:27 Decoupled.scala 249:36]
  wire  do_enq = empty ? _GEN_10 : _do_enq_T; // @[Decoupled.scala 246:18]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 246:18 Decoupled.scala 248:14]
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_resp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = 1'h0;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 245:25 Decoupled.scala 245:40 Decoupled.scala 240:16]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_resp = empty ? io_enq_bits_resp : ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_last = empty ? io_enq_bits_last : ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      if (empty) begin // @[Decoupled.scala 246:18]
        if (io_deq_ready) begin // @[Decoupled.scala 249:27]
          maybe_full <= 1'h0; // @[Decoupled.scala 249:36]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_3[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_12(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input        io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_deq_ready,
  output       io_deq_valid,
  output       io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  ram_id [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_resp [0:0]; // @[Decoupled.scala 218:16]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 249:27 Decoupled.scala 249:36]
  wire  do_enq = empty ? _GEN_8 : _do_enq_T; // @[Decoupled.scala 246:18]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 246:18 Decoupled.scala 248:14]
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_8 : _do_enq_T;
  assign ram_resp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = 1'h0;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = empty ? _GEN_8 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 245:25 Decoupled.scala 245:40 Decoupled.scala 240:16]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_resp = empty ? io_enq_bits_resp : ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      if (empty) begin // @[Decoupled.scala 246:18]
        if (io_deq_ready) begin // @[Decoupled.scala 249:27]
          maybe_full <= 1'h0; // @[Decoupled.scala 249:36]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4ToTL(
  input         clock,
  input         reset,
  output        auto_in_awready,
  input         auto_in_awvalid,
  input         auto_in_awid,
  input  [31:0] auto_in_awaddr,
  input  [7:0]  auto_in_awlen,
  input  [2:0]  auto_in_awsize,
  output        auto_in_wready,
  input         auto_in_wvalid,
  input  [63:0] auto_in_wdata,
  input  [7:0]  auto_in_wstrb,
  input         auto_in_wlast,
  input         auto_in_bready,
  output        auto_in_bvalid,
  output        auto_in_bid,
  output [1:0]  auto_in_bresp,
  output        auto_in_arready,
  input         auto_in_arvalid,
  input         auto_in_arid,
  input  [31:0] auto_in_araddr,
  input  [7:0]  auto_in_arlen,
  input  [2:0]  auto_in_arsize,
  input         auto_in_rready,
  output        auto_in_rvalid,
  output        auto_in_rid,
  output [63:0] auto_in_rdata,
  output [1:0]  auto_in_rresp,
  output        auto_in_rlast,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [2:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  deq_clock; // @[Decoupled.scala 296:21]
  wire  deq_reset; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [63:0] deq_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] deq_io_enq_bits_resp; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [63:0] deq_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] deq_io_deq_bits_resp; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_bits_last; // @[Decoupled.scala 296:21]
  wire  q_bdeq_clock; // @[Decoupled.scala 296:21]
  wire  q_bdeq_reset; // @[Decoupled.scala 296:21]
  wire  q_bdeq_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_bdeq_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  q_bdeq_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [1:0] q_bdeq_io_enq_bits_resp; // @[Decoupled.scala 296:21]
  wire  q_bdeq_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_bdeq_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  q_bdeq_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [1:0] q_bdeq_io_deq_bits_resp; // @[Decoupled.scala 296:21]
  wire [15:0] _rsize1_T = {auto_in_arlen,8'hff}; // @[Cat.scala 30:58]
  wire [22:0] _GEN_16 = {{7'd0}, _rsize1_T}; // @[Bundles.scala 31:21]
  wire [22:0] _rsize1_T_1 = _GEN_16 << auto_in_arsize; // @[Bundles.scala 31:21]
  wire [14:0] r_size_lo = _rsize1_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [15:0] _rsize_T = {r_size_lo, 1'h0}; // @[package.scala 232:35]
  wire [15:0] _rsize_T_1 = _rsize_T | 16'h1; // @[package.scala 232:40]
  wire [15:0] _rsize_T_2 = {1'h0,r_size_lo}; // @[Cat.scala 30:58]
  wire [15:0] _rsize_T_3 = ~_rsize_T_2; // @[package.scala 232:53]
  wire [15:0] _rsize_T_4 = _rsize_T_1 & _rsize_T_3; // @[package.scala 232:51]
  wire [7:0] r_size_hi = _rsize_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] r_size_lo_1 = _rsize_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  r_size_hi_1 = |r_size_hi; // @[OneHot.scala 32:14]
  wire [7:0] _rsize_T_5 = r_size_hi | r_size_lo_1; // @[OneHot.scala 32:28]
  wire [3:0] r_size_hi_2 = _rsize_T_5[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] r_size_lo_2 = _rsize_T_5[3:0]; // @[OneHot.scala 31:18]
  wire  r_size_hi_3 = |r_size_hi_2; // @[OneHot.scala 32:14]
  wire [3:0] _rsize_T_6 = r_size_hi_2 | r_size_lo_2; // @[OneHot.scala 32:28]
  wire [1:0] r_size_hi_4 = _rsize_T_6[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] r_size_lo_3 = _rsize_T_6[1:0]; // @[OneHot.scala 31:18]
  wire  r_size_hi_5 = |r_size_hi_4; // @[OneHot.scala 32:14]
  wire [1:0] _rsize_T_7 = r_size_hi_4 | r_size_lo_3; // @[OneHot.scala 32:28]
  wire  r_size_lo_4 = _rsize_T_7[1]; // @[CircuitMath.scala 30:8]
  wire [3:0] r_size = {r_size_hi_1,r_size_hi_3,r_size_hi_5,r_size_lo_4}; // @[Cat.scala 30:58]
  wire  _rok_T_1 = r_size <= 4'h6; // @[Parameters.scala 92:42]
  wire [31:0] _rok_T_4 = auto_in_araddr ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _rok_T_5 = {1'b0,$signed(_rok_T_4)}; // @[Parameters.scala 137:49]
  wire [32:0] _rok_T_7 = $signed(_rok_T_5) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _rok_T_8 = $signed(_rok_T_7) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _rok_T_9 = auto_in_araddr ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _rok_T_10 = {1'b0,$signed(_rok_T_9)}; // @[Parameters.scala 137:49]
  wire [32:0] _rok_T_12 = $signed(_rok_T_10) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _rok_T_13 = $signed(_rok_T_12) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _rok_T_14 = auto_in_araddr ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _rok_T_15 = {1'b0,$signed(_rok_T_14)}; // @[Parameters.scala 137:49]
  wire [32:0] _rok_T_17 = $signed(_rok_T_15) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _rok_T_18 = $signed(_rok_T_17) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _rok_T_19 = auto_in_araddr ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _rok_T_20 = {1'b0,$signed(_rok_T_19)}; // @[Parameters.scala 137:49]
  wire [32:0] _rok_T_22 = $signed(_rok_T_20) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _rok_T_23 = $signed(_rok_T_22) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _rok_T_24 = auto_in_araddr ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _rok_T_25 = {1'b0,$signed(_rok_T_24)}; // @[Parameters.scala 137:49]
  wire [32:0] _rok_T_27 = $signed(_rok_T_25) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _rok_T_28 = $signed(_rok_T_27) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _rok_T_32 = _rok_T_8 | _rok_T_13 | _rok_T_18 | _rok_T_23 | _rok_T_28; // @[Parameters.scala 671:42]
  wire  r_ok = _rok_T_1 & _rok_T_32; // @[Parameters.scala 670:56]
  wire [12:0] _GEN_17 = {{10'd0}, auto_in_araddr[2:0]}; // @[ToTL.scala 90:59]
  wire [12:0] _raddr_T_1 = 13'h1000 | _GEN_17; // @[ToTL.scala 90:59]
  wire [31:0] r_addr = r_ok ? auto_in_araddr : {{19'd0}, _raddr_T_1}; // @[ToTL.scala 90:23]
  reg [2:0] r_count_0; // @[ToTL.scala 91:28]
  reg [2:0] r_count_1; // @[ToTL.scala 91:28]
  wire [2:0] _GEN_1 = auto_in_arid ? r_count_1 : r_count_0; // @[ToTL.scala 95:50 ToTL.scala 95:50]
  wire [1:0] r_id_hi_lo = _GEN_1[1:0]; // @[ToTL.scala 95:50]
  wire [3:0] r_id = {auto_in_arid,r_id_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [29:0] _T_2 = 30'h7fff << r_size; // @[package.scala 234:77]
  wire [14:0] _T_4 = ~_T_2[14:0]; // @[package.scala 234:46]
  wire [1:0] a_mask_sizeOH_shiftAmount = r_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _a_mask_sizeOH_T_1 = 4'h1 << a_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] a_mask_sizeOH = _a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _a_mask_T = r_size >= 4'h3; // @[Misc.scala 205:21]
  wire  a_mask_size = a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  a_mask_bit = r_addr[2]; // @[Misc.scala 209:26]
  wire  a_mask_nbit = ~a_mask_bit; // @[Misc.scala 210:20]
  wire  a_mask_acc = _a_mask_T | a_mask_size & a_mask_nbit; // @[Misc.scala 214:29]
  wire  a_mask_acc_1 = _a_mask_T | a_mask_size & a_mask_bit; // @[Misc.scala 214:29]
  wire  a_mask_size_1 = a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  a_mask_bit_1 = r_addr[1]; // @[Misc.scala 209:26]
  wire  a_mask_nbit_1 = ~a_mask_bit_1; // @[Misc.scala 210:20]
  wire  a_mask_eq_2 = a_mask_nbit & a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_2 = a_mask_acc | a_mask_size_1 & a_mask_eq_2; // @[Misc.scala 214:29]
  wire  a_mask_eq_3 = a_mask_nbit & a_mask_bit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_3 = a_mask_acc | a_mask_size_1 & a_mask_eq_3; // @[Misc.scala 214:29]
  wire  a_mask_eq_4 = a_mask_bit & a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_4 = a_mask_acc_1 | a_mask_size_1 & a_mask_eq_4; // @[Misc.scala 214:29]
  wire  a_mask_eq_5 = a_mask_bit & a_mask_bit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_5 = a_mask_acc_1 | a_mask_size_1 & a_mask_eq_5; // @[Misc.scala 214:29]
  wire  a_mask_size_2 = a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  a_mask_bit_2 = r_addr[0]; // @[Misc.scala 209:26]
  wire  a_mask_nbit_2 = ~a_mask_bit_2; // @[Misc.scala 210:20]
  wire  a_mask_eq_6 = a_mask_eq_2 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_lo_lo_lo = a_mask_acc_2 | a_mask_size_2 & a_mask_eq_6; // @[Misc.scala 214:29]
  wire  a_mask_eq_7 = a_mask_eq_2 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_lo_lo_hi = a_mask_acc_2 | a_mask_size_2 & a_mask_eq_7; // @[Misc.scala 214:29]
  wire  a_mask_eq_8 = a_mask_eq_3 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_lo_hi_lo = a_mask_acc_3 | a_mask_size_2 & a_mask_eq_8; // @[Misc.scala 214:29]
  wire  a_mask_eq_9 = a_mask_eq_3 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_lo_hi_hi = a_mask_acc_3 | a_mask_size_2 & a_mask_eq_9; // @[Misc.scala 214:29]
  wire  a_mask_eq_10 = a_mask_eq_4 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_hi_lo_lo = a_mask_acc_4 | a_mask_size_2 & a_mask_eq_10; // @[Misc.scala 214:29]
  wire  a_mask_eq_11 = a_mask_eq_4 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_hi_lo_hi = a_mask_acc_4 | a_mask_size_2 & a_mask_eq_11; // @[Misc.scala 214:29]
  wire  a_mask_eq_12 = a_mask_eq_5 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_hi_hi_lo = a_mask_acc_5 | a_mask_size_2 & a_mask_eq_12; // @[Misc.scala 214:29]
  wire  a_mask_eq_13 = a_mask_eq_5 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_hi_hi_hi = a_mask_acc_5 | a_mask_size_2 & a_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] a_mask = {a_mask_hi_hi_hi,a_mask_hi_hi_lo,a_mask_hi_lo_hi,a_mask_hi_lo_lo,a_mask_lo_hi_hi,a_mask_lo_hi_lo,
    a_mask_lo_lo_hi,a_mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [1:0] r_sel = 2'h1 << auto_in_arid; // @[OneHot.scala 65:12]
  reg [7:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 8'h0; // @[Arbiter.scala 88:28]
  wire  w_out_valid = auto_in_awvalid & auto_in_wvalid; // @[ToTL.scala 135:34]
  wire [1:0] readys_filter_lo = {w_out_valid,auto_in_arvalid}; // @[Cat.scala 30:58]
  reg [1:0] readys_mask; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 24:30]
  wire [1:0] readys_filter_hi = readys_filter_lo & _readys_filter_T; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter = {readys_filter_hi,w_out_valid,auto_in_arvalid}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_18 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_18; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_19 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready = _GEN_19 | _readys_unready_T_4; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  wire  readys_0 = readys_readys[0]; // @[Arbiter.scala 95:86]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  out_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  wire  _T_12 = out_ready & auto_in_arvalid; // @[Decoupled.scala 40:37]
  wire [2:0] _rcount_0_T_1 = r_count_0 + 3'h1; // @[ToTL.scala 116:43]
  wire [2:0] _rcount_1_T_1 = r_count_1 + 3'h1; // @[ToTL.scala 116:43]
  wire [15:0] _wsize1_T = {auto_in_awlen,8'hff}; // @[Cat.scala 30:58]
  wire [22:0] _GEN_20 = {{7'd0}, _wsize1_T}; // @[Bundles.scala 31:21]
  wire [22:0] _wsize1_T_1 = _GEN_20 << auto_in_awsize; // @[Bundles.scala 31:21]
  wire [14:0] w_size_lo = _wsize1_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [15:0] _wsize_T = {w_size_lo, 1'h0}; // @[package.scala 232:35]
  wire [15:0] _wsize_T_1 = _wsize_T | 16'h1; // @[package.scala 232:40]
  wire [15:0] _wsize_T_2 = {1'h0,w_size_lo}; // @[Cat.scala 30:58]
  wire [15:0] _wsize_T_3 = ~_wsize_T_2; // @[package.scala 232:53]
  wire [15:0] _wsize_T_4 = _wsize_T_1 & _wsize_T_3; // @[package.scala 232:51]
  wire [7:0] w_size_hi = _wsize_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] w_size_lo_1 = _wsize_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  w_size_hi_1 = |w_size_hi; // @[OneHot.scala 32:14]
  wire [7:0] _wsize_T_5 = w_size_hi | w_size_lo_1; // @[OneHot.scala 32:28]
  wire [3:0] w_size_hi_2 = _wsize_T_5[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] w_size_lo_2 = _wsize_T_5[3:0]; // @[OneHot.scala 31:18]
  wire  w_size_hi_3 = |w_size_hi_2; // @[OneHot.scala 32:14]
  wire [3:0] _wsize_T_6 = w_size_hi_2 | w_size_lo_2; // @[OneHot.scala 32:28]
  wire [1:0] w_size_hi_4 = _wsize_T_6[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] w_size_lo_3 = _wsize_T_6[1:0]; // @[OneHot.scala 31:18]
  wire  w_size_hi_5 = |w_size_hi_4; // @[OneHot.scala 32:14]
  wire [1:0] _wsize_T_7 = w_size_hi_4 | w_size_lo_3; // @[OneHot.scala 32:28]
  wire  w_size_lo_4 = _wsize_T_7[1]; // @[CircuitMath.scala 30:8]
  wire [3:0] w_size = {w_size_hi_1,w_size_hi_3,w_size_hi_5,w_size_lo_4}; // @[Cat.scala 30:58]
  wire  _wok_T_1 = w_size <= 4'h6; // @[Parameters.scala 92:42]
  wire [31:0] _wok_T_4 = auto_in_awaddr ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _wok_T_5 = {1'b0,$signed(_wok_T_4)}; // @[Parameters.scala 137:49]
  wire [32:0] _wok_T_7 = $signed(_wok_T_5) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _wok_T_8 = $signed(_wok_T_7) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _wok_T_9 = auto_in_awaddr ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _wok_T_10 = {1'b0,$signed(_wok_T_9)}; // @[Parameters.scala 137:49]
  wire [32:0] _wok_T_12 = $signed(_wok_T_10) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _wok_T_13 = $signed(_wok_T_12) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _wok_T_14 = auto_in_awaddr ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _wok_T_15 = {1'b0,$signed(_wok_T_14)}; // @[Parameters.scala 137:49]
  wire [32:0] _wok_T_17 = $signed(_wok_T_15) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _wok_T_18 = $signed(_wok_T_17) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _wok_T_19 = auto_in_awaddr ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _wok_T_20 = {1'b0,$signed(_wok_T_19)}; // @[Parameters.scala 137:49]
  wire [32:0] _wok_T_22 = $signed(_wok_T_20) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _wok_T_23 = $signed(_wok_T_22) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _wok_T_24 = auto_in_awaddr ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _wok_T_25 = {1'b0,$signed(_wok_T_24)}; // @[Parameters.scala 137:49]
  wire [32:0] _wok_T_27 = $signed(_wok_T_25) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _wok_T_28 = $signed(_wok_T_27) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _wok_T_32 = _wok_T_8 | _wok_T_13 | _wok_T_18 | _wok_T_23 | _wok_T_28; // @[Parameters.scala 671:42]
  wire  w_ok = _wok_T_1 & _wok_T_32; // @[Parameters.scala 670:56]
  wire [12:0] _GEN_21 = {{10'd0}, auto_in_awaddr[2:0]}; // @[ToTL.scala 123:59]
  wire [12:0] _waddr_T_1 = 13'h1000 | _GEN_21; // @[ToTL.scala 123:59]
  wire [31:0] w_addr = w_ok ? auto_in_awaddr : {{19'd0}, _waddr_T_1}; // @[ToTL.scala 123:23]
  reg [2:0] w_count_0; // @[ToTL.scala 124:28]
  reg [2:0] w_count_1; // @[ToTL.scala 124:28]
  wire [2:0] _GEN_5 = auto_in_awid ? w_count_1 : w_count_0; // @[ToTL.scala 128:50 ToTL.scala 128:50]
  wire [1:0] w_id_hi_lo = _GEN_5[1:0]; // @[ToTL.scala 128:50]
  wire [3:0] w_id = {auto_in_awid,w_id_hi_lo,1'h1}; // @[Cat.scala 30:58]
  wire  _T_16 = ~auto_in_awvalid; // @[ToTL.scala 131:15]
  wire [29:0] _T_18 = 30'h7fff << w_size; // @[package.scala 234:77]
  wire [14:0] _T_20 = ~_T_18[14:0]; // @[package.scala 234:46]
  wire  readys_1 = readys_readys[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 123:31]
  wire  bundleIn_0_awready = out_1_ready & auto_in_wvalid & auto_in_wlast; // @[ToTL.scala 133:48]
  wire [1:0] w_sel = 2'h1 << auto_in_awid; // @[OneHot.scala 65:12]
  wire  _T_36 = bundleIn_0_awready & auto_in_awvalid; // @[Decoupled.scala 40:37]
  wire [2:0] _wcount_0_T_1 = w_count_0 + 3'h1; // @[ToTL.scala 152:43]
  wire [2:0] _wcount_1_T_1 = w_count_1 + 3'h1; // @[ToTL.scala 152:43]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _readys_mask_T = readys_readys & readys_filter_lo; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 244:43]
  wire  earlyWinner_0 = readys_0 & auto_in_arvalid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1 = readys_1 & w_out_valid; // @[Arbiter.scala 97:79]
  wire  _prefixOR_T = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 104:53]
  wire  _T_50 = auto_in_arvalid | w_out_valid; // @[Arbiter.scala 107:36]
  wire  _T_51 = ~(auto_in_arvalid | w_out_valid); // @[Arbiter.scala 107:15]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & auto_in_arvalid | state_1 & w_out_valid; // @[Mux.scala 27:72]
  wire  sink_ACancel_earlyValid = idle ? _T_50 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 50:33]
  wire [7:0] _GEN_22 = {{7'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [7:0] _beatsLeft_T_4 = beatsLeft - _GEN_22; // @[Arbiter.scala 113:52]
  wire [7:0] _T_70 = muxStateEarly_0 ? a_mask : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_71 = muxStateEarly_1 ? auto_in_wstrb : 8'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_73 = muxStateEarly_0 ? r_addr : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_74 = muxStateEarly_1 ? w_addr : 32'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_76 = muxStateEarly_0 ? r_id : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_77 = muxStateEarly_1 ? w_id : 4'h0; // @[Mux.scala 27:72]
  wire [2:0] a_size = r_size[2:0]; // @[Edges.scala 447:17 Edges.scala 450:15]
  wire [2:0] _T_79 = muxStateEarly_0 ? a_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] a_1_size = w_size[2:0]; // @[Edges.scala 483:17 Edges.scala 486:15]
  wire [2:0] _T_80 = muxStateEarly_1 ? a_1_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_85 = muxStateEarly_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_86 = muxStateEarly_1 ? 3'h1 : 3'h0; // @[Mux.scala 27:72]
  wire  d_hasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  ok_rready = deq_io_enq_ready; // @[ToTL.scala 158:23 Decoupled.scala 299:17]
  wire  ok_bready = q_bdeq_io_enq_ready; // @[ToTL.scala 157:23 Decoupled.scala 299:17]
  wire  bundleOut_0_d_ready = d_hasData ? ok_rready : ok_bready; // @[ToTL.scala 164:25]
  wire  _d_last_T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_last_beats1_decode_T_1 = 13'h3f << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_last_beats1_decode_T_3 = ~_d_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_last_beats1_decode = _d_last_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire [2:0] d_last_beats1 = d_hasData ? d_last_beats1_decode : 3'h0; // @[Edges.scala 220:14]
  reg [2:0] d_last_counter; // @[Edges.scala 228:27]
  wire [2:0] d_last_counter1 = d_last_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_last_first = d_last_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] b_count_0; // @[ToTL.scala 186:28]
  reg [2:0] b_count_1; // @[ToTL.scala 186:28]
  wire  q_bid = q_bdeq_io_deq_bits_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire [2:0] _GEN_11 = q_bid ? b_count_1 : b_count_0; // @[ToTL.scala 187:43 ToTL.scala 187:43]
  wire [2:0] _GEN_13 = q_bid ? w_count_1 : w_count_0; // @[ToTL.scala 187:43 ToTL.scala 187:43]
  wire  b_allow = _GEN_11 != _GEN_13; // @[ToTL.scala 187:43]
  wire [1:0] b_sel = 2'h1 << q_bid; // @[OneHot.scala 65:12]
  wire  q_bvalid = q_bdeq_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  bundleIn_0_bvalid = q_bvalid & b_allow; // @[ToTL.scala 195:31]
  wire  _T_90 = auto_in_bready & bundleIn_0_bvalid; // @[Decoupled.scala 40:37]
  wire [2:0] _bcount_0_T_1 = b_count_0 + 3'h1; // @[ToTL.scala 191:42]
  wire [2:0] _bcount_1_T_1 = b_count_1 + 3'h1; // @[ToTL.scala 191:42]
  Queue_11 deq ( // @[Decoupled.scala 296:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_id(deq_io_enq_bits_id),
    .io_enq_bits_data(deq_io_enq_bits_data),
    .io_enq_bits_resp(deq_io_enq_bits_resp),
    .io_enq_bits_last(deq_io_enq_bits_last),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_id(deq_io_deq_bits_id),
    .io_deq_bits_data(deq_io_deq_bits_data),
    .io_deq_bits_resp(deq_io_deq_bits_resp),
    .io_deq_bits_last(deq_io_deq_bits_last)
  );
  Queue_12 q_bdeq ( // @[Decoupled.scala 296:21]
    .clock(q_bdeq_clock),
    .reset(q_bdeq_reset),
    .io_enq_ready(q_bdeq_io_enq_ready),
    .io_enq_valid(q_bdeq_io_enq_valid),
    .io_enq_bits_id(q_bdeq_io_enq_bits_id),
    .io_enq_bits_resp(q_bdeq_io_enq_bits_resp),
    .io_deq_ready(q_bdeq_io_deq_ready),
    .io_deq_valid(q_bdeq_io_deq_valid),
    .io_deq_bits_id(q_bdeq_io_deq_bits_id),
    .io_deq_bits_resp(q_bdeq_io_deq_bits_resp)
  );
  assign auto_in_awready = out_1_ready & auto_in_wvalid & auto_in_wlast; // @[ToTL.scala 133:48]
  assign auto_in_wready = out_1_ready & auto_in_awvalid; // @[ToTL.scala 134:34]
  assign auto_in_bvalid = q_bvalid & b_allow; // @[ToTL.scala 195:31]
  assign auto_in_bid = q_bdeq_io_deq_bits_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_in_bresp = q_bdeq_io_deq_bits_resp; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_in_arready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  assign auto_in_rvalid = deq_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  assign auto_in_rid = deq_io_deq_bits_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_in_rdata = deq_io_deq_bits_data; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_in_rresp = deq_io_deq_bits_resp; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_in_rlast = deq_io_deq_bits_last; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_a_valid = idle ? _T_50 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_out_a_bits_opcode = _T_85 | _T_86; // @[Mux.scala 27:72]
  assign auto_out_a_bits_size = _T_79 | _T_80; // @[Mux.scala 27:72]
  assign auto_out_a_bits_source = _T_76 | _T_77; // @[Mux.scala 27:72]
  assign auto_out_a_bits_address = _T_73 | _T_74; // @[Mux.scala 27:72]
  assign auto_out_a_bits_mask = _T_70 | _T_71; // @[Mux.scala 27:72]
  assign auto_out_a_bits_data = muxStateEarly_1 ? auto_in_wdata : 64'h0; // @[Mux.scala 27:72]
  assign auto_out_d_ready = d_hasData ? ok_rready : ok_bready; // @[ToTL.scala 164:25]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = auto_out_d_valid & d_hasData; // @[ToTL.scala 165:33]
  assign deq_io_enq_bits_id = auto_out_d_bits_source[3]; // @[ToTL.scala 168:43]
  assign deq_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign deq_io_enq_bits_resp = auto_out_d_bits_denied | auto_out_d_bits_corrupt ? 2'h2 : 2'h0; // @[ToTL.scala 160:23]
  assign deq_io_enq_bits_last = d_last_counter == 3'h1 | d_last_beats1 == 3'h0; // @[Edges.scala 231:37]
  assign deq_io_deq_ready = auto_in_rready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign q_bdeq_clock = clock;
  assign q_bdeq_reset = reset;
  assign q_bdeq_io_enq_valid = auto_out_d_valid & ~d_hasData; // @[ToTL.scala 166:33]
  assign q_bdeq_io_enq_bits_id = auto_out_d_bits_source[3]; // @[ToTL.scala 177:43]
  assign q_bdeq_io_enq_bits_resp = auto_out_d_bits_denied | auto_out_d_bits_corrupt ? 2'h2 : 2'h0; // @[ToTL.scala 160:23]
  assign q_bdeq_io_deq_ready = auto_in_bready & b_allow; // @[ToTL.scala 196:31]
  always @(posedge clock) begin
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_0 <= 3'h0; // @[ToTL.scala 91:28]
    end else if (_T_12 & r_sel[0]) begin // @[ToTL.scala 116:34]
      r_count_0 <= _rcount_0_T_1; // @[ToTL.scala 116:38]
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_1 <= 3'h0; // @[ToTL.scala 91:28]
    end else if (_T_12 & r_sel[1]) begin // @[ToTL.scala 116:34]
      r_count_1 <= _rcount_1_T_1; // @[ToTL.scala 116:38]
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 8'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin // @[Arbiter.scala 113:23]
      if (earlyWinner_1) begin // @[Arbiter.scala 111:73]
        beatsLeft <= auto_in_awlen;
      end else begin
        beatsLeft <= 8'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch & |readys_filter_lo) begin // @[Arbiter.scala 27:32]
      readys_mask <= _readys_mask_T_3; // @[Arbiter.scala 28:12]
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin // @[Arbiter.scala 117:30]
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_0 <= 3'h0; // @[ToTL.scala 124:28]
    end else if (_T_36 & w_sel[0]) begin // @[ToTL.scala 152:34]
      w_count_0 <= _wcount_0_T_1; // @[ToTL.scala 152:38]
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_1 <= 3'h0; // @[ToTL.scala 124:28]
    end else if (_T_36 & w_sel[1]) begin // @[ToTL.scala 152:34]
      w_count_1 <= _wcount_1_T_1; // @[ToTL.scala 152:38]
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin // @[Arbiter.scala 117:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_last_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_last_T) begin // @[Edges.scala 234:17]
      if (d_last_first) begin // @[Edges.scala 235:21]
        if (d_hasData) begin // @[Edges.scala 220:14]
          d_last_counter <= d_last_beats1_decode;
        end else begin
          d_last_counter <= 3'h0;
        end
      end else begin
        d_last_counter <= d_last_counter1;
      end
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_0 <= 3'h0; // @[ToTL.scala 186:28]
    end else if (_T_90 & b_sel[0]) begin // @[ToTL.scala 191:33]
      b_count_0 <= _bcount_0_T_1; // @[ToTL.scala 191:37]
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_1 <= 3'h0; // @[ToTL.scala 186:28]
    end else if (_T_90 & b_sel[1]) begin // @[ToTL.scala 191:33]
      b_count_1 <= _bcount_1_T_1; // @[ToTL.scala 191:37]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~auto_in_arvalid | r_size_lo == _T_4 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:98 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n"
            ); // @[ToTL.scala 98:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_in_arvalid | r_size_lo == _T_4 | reset)) begin
          $fatal; // @[ToTL.scala 98:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~auto_in_awvalid | w_size_lo == _T_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:131 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n"
            ); // @[ToTL.scala 131:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_in_awvalid | w_size_lo == _T_20 | reset)) begin
          $fatal; // @[ToTL.scala 131:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_16 | auto_in_awlen == 8'h0 | auto_in_awsize == 3'h3 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:132 assert (!in.aw.valid || in.aw.bits.len === UInt(0) || in.aw.bits.size === UInt(log2Ceil(beatBytes))) // because aligned\n"
            ); // @[ToTL.scala 132:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_16 | auto_in_awlen == 8'h0 | auto_in_awsize == 3'h3 | reset)) begin
          $fatal; // @[ToTL.scala 132:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(auto_in_arvalid | w_out_valid) | _prefixOR_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(auto_in_arvalid | w_out_valid) | _prefixOR_T | reset)) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_51 | _T_50 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_51 | _T_50 | reset)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_count_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  r_count_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  beatsLeft = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  readys_mask = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  state_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  w_count_0 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  w_count_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  state_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  d_last_counter = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  b_count_0 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  b_count_1 = _RAND_10[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueCompatibility(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_extra_id,
  input        io_enq_bits_real_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_extra_id,
  output       io_deq_bits_real_last
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_extra_id [0:3]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [1:0] ram_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_extra_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [1:0] ram_extra_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_real_last [0:3]; // @[Decoupled.scala 218:16]
  wire  ram_real_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [1:0] ram_real_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_real_last_MPORT_data; // @[Decoupled.scala 218:16]
  wire [1:0] ram_real_last_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_real_last_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_real_last_MPORT_en; // @[Decoupled.scala 218:16]
  reg [1:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 76:24]
  wire  _GEN_10 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 249:27 Decoupled.scala 249:36]
  wire  do_enq = empty ? _GEN_10 : _do_enq_T; // @[Decoupled.scala 246:18]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 76:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 246:18 Decoupled.scala 248:14]
  assign ram_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_extra_id_MPORT_data = io_enq_bits_extra_id;
  assign ram_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_extra_id_MPORT_mask = 1'h1;
  assign ram_extra_id_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_real_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_real_last_io_deq_bits_MPORT_data = ram_real_last[ram_real_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_real_last_MPORT_data = io_enq_bits_real_last;
  assign ram_real_last_MPORT_addr = enq_ptr_value;
  assign ram_real_last_MPORT_mask = 1'h1;
  assign ram_real_last_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 245:25 Decoupled.scala 245:40 Decoupled.scala 240:16]
  assign io_deq_bits_extra_id = empty ? io_enq_bits_extra_id : ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_real_last = empty ? io_enq_bits_real_last : ram_real_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_extra_id_MPORT_en & ram_extra_id_MPORT_mask) begin
      ram_extra_id[ram_extra_id_MPORT_addr] <= ram_extra_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_real_last_MPORT_en & ram_real_last_MPORT_mask) begin
      ram_real_last[ram_real_last_MPORT_addr] <= ram_real_last_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      if (empty) begin // @[Decoupled.scala 246:18]
        if (io_deq_ready) begin // @[Decoupled.scala 249:27]
          maybe_full <= 1'h0; // @[Decoupled.scala 249:36]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_extra_id[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_real_last[initvar] = _RAND_1[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4UserYanker(
  input         clock,
  input         reset,
  output        auto_in_awready,
  input         auto_in_awvalid,
  input         auto_in_awid,
  input  [31:0] auto_in_awaddr,
  input  [7:0]  auto_in_awlen,
  input  [2:0]  auto_in_awsize,
  input  [2:0]  auto_in_awecho_extra_id,
  input         auto_in_awecho_real_last,
  output        auto_in_wready,
  input         auto_in_wvalid,
  input  [63:0] auto_in_wdata,
  input  [7:0]  auto_in_wstrb,
  input         auto_in_wlast,
  input         auto_in_bready,
  output        auto_in_bvalid,
  output        auto_in_bid,
  output [1:0]  auto_in_bresp,
  output [2:0]  auto_in_becho_extra_id,
  output        auto_in_becho_real_last,
  output        auto_in_arready,
  input         auto_in_arvalid,
  input         auto_in_arid,
  input  [31:0] auto_in_araddr,
  input  [7:0]  auto_in_arlen,
  input  [2:0]  auto_in_arsize,
  input  [2:0]  auto_in_arecho_extra_id,
  input         auto_in_arecho_real_last,
  input         auto_in_rready,
  output        auto_in_rvalid,
  output        auto_in_rid,
  output [63:0] auto_in_rdata,
  output [1:0]  auto_in_rresp,
  output [2:0]  auto_in_recho_extra_id,
  output        auto_in_recho_real_last,
  output        auto_in_rlast,
  input         auto_out_awready,
  output        auto_out_awvalid,
  output        auto_out_awid,
  output [31:0] auto_out_awaddr,
  output [7:0]  auto_out_awlen,
  output [2:0]  auto_out_awsize,
  input         auto_out_wready,
  output        auto_out_wvalid,
  output [63:0] auto_out_wdata,
  output [7:0]  auto_out_wstrb,
  output        auto_out_wlast,
  output        auto_out_bready,
  input         auto_out_bvalid,
  input         auto_out_bid,
  input  [1:0]  auto_out_bresp,
  input         auto_out_arready,
  output        auto_out_arvalid,
  output        auto_out_arid,
  output [31:0] auto_out_araddr,
  output [7:0]  auto_out_arlen,
  output [2:0]  auto_out_arsize,
  output        auto_out_rready,
  input         auto_out_rvalid,
  input         auto_out_rid,
  input  [63:0] auto_out_rdata,
  input  [1:0]  auto_out_rresp,
  input         auto_out_rlast
);
  wire  QueueCompatibility_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [2:0] QueueCompatibility_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [2:0] QueueCompatibility_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [2:0] QueueCompatibility_1_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [2:0] QueueCompatibility_1_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [2:0] QueueCompatibility_2_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [2:0] QueueCompatibility_2_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [2:0] QueueCompatibility_3_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [2:0] QueueCompatibility_3_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  _arready_WIRE_0 = QueueCompatibility_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _arready_WIRE_1 = QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_1 = auto_in_arid ? _arready_WIRE_1 : _arready_WIRE_0; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _rvalid_WIRE_0 = QueueCompatibility_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _rvalid_WIRE_1 = QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_3 = auto_out_rid ? _rvalid_WIRE_1 : _rvalid_WIRE_0; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rWIRE_0_real_last = QueueCompatibility_io_deq_bits_real_last; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _rWIRE_1_real_last = QueueCompatibility_1_io_deq_bits_real_last; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [2:0] _rWIRE_0_extra_id = QueueCompatibility_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [2:0] _rWIRE_1_extra_id = QueueCompatibility_1_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [1:0] _arsel_T = 2'h1 << auto_in_arid; // @[OneHot.scala 65:12]
  wire  arsel_0 = _arsel_T[0]; // @[UserYanker.scala 67:55]
  wire  arsel_1 = _arsel_T[1]; // @[UserYanker.scala 67:55]
  wire [1:0] _rsel_T = 2'h1 << auto_out_rid; // @[OneHot.scala 65:12]
  wire  rsel_0 = _rsel_T[0]; // @[UserYanker.scala 68:55]
  wire  rsel_1 = _rsel_T[1]; // @[UserYanker.scala 68:55]
  wire  _awready_WIRE_0 = QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _awready_WIRE_1 = QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_9 = auto_in_awid ? _awready_WIRE_1 : _awready_WIRE_0; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _bvalid_WIRE_0 = QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _bvalid_WIRE_1 = QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_11 = auto_out_bid ? _bvalid_WIRE_1 : _bvalid_WIRE_0; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bWIRE_0_real_last = QueueCompatibility_2_io_deq_bits_real_last; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _bWIRE_1_real_last = QueueCompatibility_3_io_deq_bits_real_last; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [2:0] _bWIRE_0_extra_id = QueueCompatibility_2_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [2:0] _bWIRE_1_extra_id = QueueCompatibility_3_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [1:0] _awsel_T = 2'h1 << auto_in_awid; // @[OneHot.scala 65:12]
  wire  awsel_0 = _awsel_T[0]; // @[UserYanker.scala 88:55]
  wire  awsel_1 = _awsel_T[1]; // @[UserYanker.scala 88:55]
  wire [1:0] _bsel_T = 2'h1 << auto_out_bid; // @[OneHot.scala 65:12]
  wire  bsel_0 = _bsel_T[0]; // @[UserYanker.scala 89:55]
  wire  bsel_1 = _bsel_T[1]; // @[UserYanker.scala 89:55]
  QueueCompatibility QueueCompatibility ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_clock),
    .reset(QueueCompatibility_reset),
    .io_enq_ready(QueueCompatibility_io_enq_ready),
    .io_enq_valid(QueueCompatibility_io_enq_valid),
    .io_enq_bits_extra_id(QueueCompatibility_io_enq_bits_extra_id),
    .io_enq_bits_real_last(QueueCompatibility_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_io_deq_ready),
    .io_deq_valid(QueueCompatibility_io_deq_valid),
    .io_deq_bits_extra_id(QueueCompatibility_io_deq_bits_extra_id),
    .io_deq_bits_real_last(QueueCompatibility_io_deq_bits_real_last)
  );
  QueueCompatibility QueueCompatibility_1 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_1_clock),
    .reset(QueueCompatibility_1_reset),
    .io_enq_ready(QueueCompatibility_1_io_enq_ready),
    .io_enq_valid(QueueCompatibility_1_io_enq_valid),
    .io_enq_bits_extra_id(QueueCompatibility_1_io_enq_bits_extra_id),
    .io_enq_bits_real_last(QueueCompatibility_1_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_1_io_deq_ready),
    .io_deq_valid(QueueCompatibility_1_io_deq_valid),
    .io_deq_bits_extra_id(QueueCompatibility_1_io_deq_bits_extra_id),
    .io_deq_bits_real_last(QueueCompatibility_1_io_deq_bits_real_last)
  );
  QueueCompatibility QueueCompatibility_2 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_2_clock),
    .reset(QueueCompatibility_2_reset),
    .io_enq_ready(QueueCompatibility_2_io_enq_ready),
    .io_enq_valid(QueueCompatibility_2_io_enq_valid),
    .io_enq_bits_extra_id(QueueCompatibility_2_io_enq_bits_extra_id),
    .io_enq_bits_real_last(QueueCompatibility_2_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_2_io_deq_ready),
    .io_deq_valid(QueueCompatibility_2_io_deq_valid),
    .io_deq_bits_extra_id(QueueCompatibility_2_io_deq_bits_extra_id),
    .io_deq_bits_real_last(QueueCompatibility_2_io_deq_bits_real_last)
  );
  QueueCompatibility QueueCompatibility_3 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_3_clock),
    .reset(QueueCompatibility_3_reset),
    .io_enq_ready(QueueCompatibility_3_io_enq_ready),
    .io_enq_valid(QueueCompatibility_3_io_enq_valid),
    .io_enq_bits_extra_id(QueueCompatibility_3_io_enq_bits_extra_id),
    .io_enq_bits_real_last(QueueCompatibility_3_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_3_io_deq_ready),
    .io_deq_valid(QueueCompatibility_3_io_deq_valid),
    .io_deq_bits_extra_id(QueueCompatibility_3_io_deq_bits_extra_id),
    .io_deq_bits_real_last(QueueCompatibility_3_io_deq_bits_real_last)
  );
  assign auto_in_awready = auto_out_awready & _GEN_9; // @[UserYanker.scala 77:36]
  assign auto_in_wready = auto_out_wready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bvalid = auto_out_bvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bid = auto_out_bid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bresp = auto_out_bresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_becho_extra_id = auto_out_bid ? _bWIRE_1_extra_id : _bWIRE_0_extra_id; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_becho_real_last = auto_out_bid ? _bWIRE_1_real_last : _bWIRE_0_real_last; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_arready = auto_out_arready & _GEN_1; // @[UserYanker.scala 56:36]
  assign auto_in_rvalid = auto_out_rvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rid = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rdata = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rresp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_recho_extra_id = auto_out_rid ? _rWIRE_1_extra_id : _rWIRE_0_extra_id; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_recho_real_last = auto_out_rid ? _rWIRE_1_real_last : _rWIRE_0_real_last; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_rlast = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_awvalid = auto_in_awvalid & _GEN_9; // @[UserYanker.scala 78:36]
  assign auto_out_awid = auto_in_awid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awaddr = auto_in_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awlen = auto_in_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awsize = auto_in_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wvalid = auto_in_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wdata = auto_in_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wstrb = auto_in_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wlast = auto_in_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_bready = auto_in_bready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arvalid = auto_in_arvalid & _GEN_1; // @[UserYanker.scala 57:36]
  assign auto_out_arid = auto_in_arid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_araddr = auto_in_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arlen = auto_in_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arsize = auto_in_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_rready = auto_in_rready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_clock = clock;
  assign QueueCompatibility_reset = reset;
  assign QueueCompatibility_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_0; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_enq_bits_real_last = auto_in_arecho_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_0 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_1_clock = clock;
  assign QueueCompatibility_1_reset = reset;
  assign QueueCompatibility_1_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_1; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_1_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_enq_bits_real_last = auto_in_arecho_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_1 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_2_clock = clock;
  assign QueueCompatibility_2_reset = reset;
  assign QueueCompatibility_2_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_0; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_2_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_enq_bits_real_last = auto_in_awecho_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_0; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_3_clock = clock;
  assign QueueCompatibility_3_reset = reset;
  assign QueueCompatibility_3_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_1; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_3_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_enq_bits_real_last = auto_in_awecho_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_1; // @[UserYanker.scala 91:53]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~auto_out_rvalid | _GEN_3 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:63 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 63:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_rvalid | _GEN_3 | reset)) begin
          $fatal; // @[UserYanker.scala 63:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~auto_out_bvalid | _GEN_11 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:84 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 84:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_bvalid | _GEN_11 | reset)) begin
          $fatal; // @[UserYanker.scala 84:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_13(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input  [2:0]  io_enq_bits_echo_extra_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [2:0]  io_deq_bits_echo_extra_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  ram_id [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_len [0:0]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_burst [0:0]; // @[Decoupled.scala 218:16]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_echo_extra_id [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_echo_extra_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_echo_extra_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_echo_extra_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_16 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 249:27 Decoupled.scala 249:36]
  wire  do_enq = empty ? _GEN_16 : _do_enq_T; // @[Decoupled.scala 246:18]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 246:18 Decoupled.scala 248:14]
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_16 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_16 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_16 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_16 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_16 : _do_enq_T;
  assign ram_echo_extra_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_extra_id_io_deq_bits_MPORT_data = ram_echo_extra_id[ram_echo_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_echo_extra_id_MPORT_data = io_enq_bits_echo_extra_id;
  assign ram_echo_extra_id_MPORT_addr = 1'h0;
  assign ram_echo_extra_id_MPORT_mask = 1'h1;
  assign ram_echo_extra_id_MPORT_en = empty ? _GEN_16 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 245:25 Decoupled.scala 245:40 Decoupled.scala 240:16]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_burst = empty ? io_enq_bits_burst : ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_echo_extra_id = empty ? io_enq_bits_echo_extra_id : ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_echo_extra_id_MPORT_en & ram_echo_extra_id_MPORT_mask) begin
      ram_echo_extra_id[ram_echo_extra_id_MPORT_addr] <= ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      if (empty) begin // @[Decoupled.scala 246:18]
        if (io_deq_ready) begin // @[Decoupled.scala 249:27]
          maybe_full <= 1'h0; // @[Decoupled.scala 249:36]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_echo_extra_id[initvar] = _RAND_5[2:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_15(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_strb,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_strb,
  output        io_deq_bits_last
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_strb [0:0]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_strb_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_strb_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_strb_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_strb_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_strb_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_last [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_9 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 249:27 Decoupled.scala 249:36]
  wire  do_enq = empty ? _GEN_9 : _do_enq_T; // @[Decoupled.scala 246:18]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 246:18 Decoupled.scala 248:14]
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_9 : _do_enq_T;
  assign ram_strb_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = 1'h0;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = empty ? _GEN_9 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_9 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 245:25 Decoupled.scala 245:40 Decoupled.scala 240:16]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_strb = empty ? io_enq_bits_strb : ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_last = empty ? io_enq_bits_last : ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      if (empty) begin // @[Decoupled.scala 246:18]
        if (io_deq_ready) begin // @[Decoupled.scala 249:27]
          maybe_full <= 1'h0; // @[Decoupled.scala 249:36]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Fragmenter(
  input         clock,
  input         reset,
  output        auto_in_awready,
  input         auto_in_awvalid,
  input         auto_in_awid,
  input  [31:0] auto_in_awaddr,
  input  [7:0]  auto_in_awlen,
  input  [2:0]  auto_in_awsize,
  input  [1:0]  auto_in_awburst,
  input  [2:0]  auto_in_awecho_extra_id,
  output        auto_in_wready,
  input         auto_in_wvalid,
  input  [63:0] auto_in_wdata,
  input  [7:0]  auto_in_wstrb,
  input         auto_in_wlast,
  input         auto_in_bready,
  output        auto_in_bvalid,
  output        auto_in_bid,
  output [1:0]  auto_in_bresp,
  output [2:0]  auto_in_becho_extra_id,
  output        auto_in_arready,
  input         auto_in_arvalid,
  input         auto_in_arid,
  input  [31:0] auto_in_araddr,
  input  [7:0]  auto_in_arlen,
  input  [2:0]  auto_in_arsize,
  input  [1:0]  auto_in_arburst,
  input  [2:0]  auto_in_arecho_extra_id,
  input         auto_in_rready,
  output        auto_in_rvalid,
  output        auto_in_rid,
  output [63:0] auto_in_rdata,
  output [1:0]  auto_in_rresp,
  output [2:0]  auto_in_recho_extra_id,
  output        auto_in_rlast,
  input         auto_out_awready,
  output        auto_out_awvalid,
  output        auto_out_awid,
  output [31:0] auto_out_awaddr,
  output [7:0]  auto_out_awlen,
  output [2:0]  auto_out_awsize,
  output [2:0]  auto_out_awecho_extra_id,
  output        auto_out_awecho_real_last,
  input         auto_out_wready,
  output        auto_out_wvalid,
  output [63:0] auto_out_wdata,
  output [7:0]  auto_out_wstrb,
  output        auto_out_wlast,
  output        auto_out_bready,
  input         auto_out_bvalid,
  input         auto_out_bid,
  input  [1:0]  auto_out_bresp,
  input  [2:0]  auto_out_becho_extra_id,
  input         auto_out_becho_real_last,
  input         auto_out_arready,
  output        auto_out_arvalid,
  output        auto_out_arid,
  output [31:0] auto_out_araddr,
  output [7:0]  auto_out_arlen,
  output [2:0]  auto_out_arsize,
  output [2:0]  auto_out_arecho_extra_id,
  output        auto_out_arecho_real_last,
  output        auto_out_rready,
  input         auto_out_rvalid,
  input         auto_out_rid,
  input  [63:0] auto_out_rdata,
  input  [1:0]  auto_out_rresp,
  input  [2:0]  auto_out_recho_extra_id,
  input         auto_out_recho_real_last,
  input         auto_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  deq_clock; // @[Decoupled.scala 296:21]
  wire  deq_reset; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [31:0] deq_io_enq_bits_addr; // @[Decoupled.scala 296:21]
  wire [7:0] deq_io_enq_bits_len; // @[Decoupled.scala 296:21]
  wire [2:0] deq_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] deq_io_enq_bits_burst; // @[Decoupled.scala 296:21]
  wire [2:0] deq_io_enq_bits_echo_extra_id; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [31:0] deq_io_deq_bits_addr; // @[Decoupled.scala 296:21]
  wire [7:0] deq_io_deq_bits_len; // @[Decoupled.scala 296:21]
  wire [2:0] deq_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] deq_io_deq_bits_burst; // @[Decoupled.scala 296:21]
  wire [2:0] deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 296:21]
  wire  deq_1_clock; // @[Decoupled.scala 296:21]
  wire  deq_1_reset; // @[Decoupled.scala 296:21]
  wire  deq_1_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  deq_1_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  deq_1_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [31:0] deq_1_io_enq_bits_addr; // @[Decoupled.scala 296:21]
  wire [7:0] deq_1_io_enq_bits_len; // @[Decoupled.scala 296:21]
  wire [2:0] deq_1_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] deq_1_io_enq_bits_burst; // @[Decoupled.scala 296:21]
  wire [2:0] deq_1_io_enq_bits_echo_extra_id; // @[Decoupled.scala 296:21]
  wire  deq_1_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  deq_1_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  deq_1_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [31:0] deq_1_io_deq_bits_addr; // @[Decoupled.scala 296:21]
  wire [7:0] deq_1_io_deq_bits_len; // @[Decoupled.scala 296:21]
  wire [2:0] deq_1_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] deq_1_io_deq_bits_burst; // @[Decoupled.scala 296:21]
  wire [2:0] deq_1_io_deq_bits_echo_extra_id; // @[Decoupled.scala 296:21]
  wire  in_wdeq_clock; // @[Decoupled.scala 296:21]
  wire  in_wdeq_reset; // @[Decoupled.scala 296:21]
  wire  in_wdeq_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  in_wdeq_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] in_wdeq_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [7:0] in_wdeq_io_enq_bits_strb; // @[Decoupled.scala 296:21]
  wire  in_wdeq_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  in_wdeq_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  in_wdeq_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] in_wdeq_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [7:0] in_wdeq_io_deq_bits_strb; // @[Decoupled.scala 296:21]
  wire  in_wdeq_io_deq_bits_last; // @[Decoupled.scala 296:21]
  reg  busy; // @[Fragmenter.scala 60:29]
  reg [31:0] r_addr; // @[Fragmenter.scala 61:25]
  reg [7:0] r_len; // @[Fragmenter.scala 62:25]
  wire [7:0] irr_bits_len = deq_io_deq_bits_len; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire [7:0] len = busy ? r_len : irr_bits_len; // @[Fragmenter.scala 64:23]
  wire [31:0] irr_bits_addr = deq_io_deq_bits_addr; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire [31:0] addr = busy ? r_addr : irr_bits_addr; // @[Fragmenter.scala 65:23]
  wire [7:0] alignment = addr[10:3]; // @[Fragmenter.scala 69:29]
  wire [7:0] _GEN_16 = {{1'd0}, len[7:1]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_1 = len | _GEN_16; // @[package.scala 253:43]
  wire [7:0] _GEN_17 = {{2'd0}, _fillLow_T_1[7:2]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_3 = _fillLow_T_1 | _GEN_17; // @[package.scala 253:43]
  wire [7:0] _GEN_18 = {{4'd0}, _fillLow_T_3[7:4]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_5 = _fillLow_T_3 | _GEN_18; // @[package.scala 253:43]
  wire [6:0] fillLow = _fillLow_T_5[7:1]; // @[Fragmenter.scala 85:37]
  wire [7:0] _wipeHigh_T = ~len; // @[Fragmenter.scala 86:32]
  wire [8:0] _wipeHigh_T_1 = {_wipeHigh_T, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_3 = _wipeHigh_T | _wipeHigh_T_1[7:0]; // @[package.scala 244:43]
  wire [9:0] _wipeHigh_T_4 = {_wipeHigh_T_3, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_6 = _wipeHigh_T_3 | _wipeHigh_T_4[7:0]; // @[package.scala 244:43]
  wire [11:0] _wipeHigh_T_7 = {_wipeHigh_T_6, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_9 = _wipeHigh_T_6 | _wipeHigh_T_7[7:0]; // @[package.scala 244:43]
  wire [7:0] wipeHigh = ~_wipeHigh_T_9; // @[Fragmenter.scala 86:24]
  wire [7:0] _GEN_19 = {{1'd0}, fillLow}; // @[Fragmenter.scala 87:32]
  wire [7:0] remain1 = _GEN_19 | wipeHigh; // @[Fragmenter.scala 87:32]
  wire [8:0] _align1_T = {alignment, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_2 = alignment | _align1_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _align1_T_3 = {_align1_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_5 = _align1_T_2 | _align1_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _align1_T_6 = {_align1_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_8 = _align1_T_5 | _align1_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] align1 = ~_align1_T_8; // @[Fragmenter.scala 88:24]
  wire [7:0] _maxSupported1_T = remain1 & align1; // @[Fragmenter.scala 89:37]
  wire [7:0] maxSupported1 = _maxSupported1_T & 8'h7; // @[Fragmenter.scala 89:46]
  wire [1:0] irr_bits_burst = deq_io_deq_bits_burst; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  fixed = irr_bits_burst == 2'h0; // @[Fragmenter.scala 92:34]
  wire [2:0] irr_bits_size = deq_io_deq_bits_size; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  narrow = irr_bits_size != 3'h3; // @[Fragmenter.scala 93:34]
  wire  bad = fixed | narrow; // @[Fragmenter.scala 94:25]
  wire [7:0] beats_lo = bad ? 8'h0 : maxSupported1; // @[Fragmenter.scala 97:25]
  wire [8:0] _beats_T = {beats_lo, 1'h0}; // @[package.scala 232:35]
  wire [8:0] _beats_T_1 = _beats_T | 9'h1; // @[package.scala 232:40]
  wire [8:0] _beats_T_2 = {1'h0,beats_lo}; // @[Cat.scala 30:58]
  wire [8:0] _beats_T_3 = ~_beats_T_2; // @[package.scala 232:53]
  wire [8:0] beats = _beats_T_1 & _beats_T_3; // @[package.scala 232:51]
  wire [15:0] _GEN_20 = {{7'd0}, beats}; // @[Fragmenter.scala 100:38]
  wire [15:0] _inc_addr_T = _GEN_20 << irr_bits_size; // @[Fragmenter.scala 100:38]
  wire [31:0] _GEN_21 = {{16'd0}, _inc_addr_T}; // @[Fragmenter.scala 100:29]
  wire [31:0] inc_addr = addr + _GEN_21; // @[Fragmenter.scala 100:29]
  wire [15:0] _wrapMask_T = {irr_bits_len,8'hff}; // @[Cat.scala 30:58]
  wire [22:0] _GEN_22 = {{7'd0}, _wrapMask_T}; // @[Bundles.scala 31:21]
  wire [22:0] _wrapMask_T_1 = _GEN_22 << irr_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] wrapMask = _wrapMask_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [31:0] _GEN_23 = {{17'd0}, wrapMask}; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T = inc_addr & _GEN_23; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_1 = ~irr_bits_addr; // @[Fragmenter.scala 104:49]
  wire [31:0] _mux_addr_T_2 = _mux_addr_T_1 | _GEN_23; // @[Fragmenter.scala 104:62]
  wire [31:0] _mux_addr_T_3 = ~_mux_addr_T_2; // @[Fragmenter.scala 104:47]
  wire [31:0] _mux_addr_T_4 = _mux_addr_T | _mux_addr_T_3; // @[Fragmenter.scala 104:45]
  wire  ar_last = beats_lo == len; // @[Fragmenter.scala 110:27]
  wire [31:0] _out_bits_addr_T = ~addr; // @[Fragmenter.scala 122:28]
  wire [9:0] _out_bits_addr_T_2 = 10'h7 << irr_bits_size; // @[package.scala 234:77]
  wire [2:0] _out_bits_addr_T_4 = ~_out_bits_addr_T_2[2:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_25 = {{29'd0}, _out_bits_addr_T_4}; // @[Fragmenter.scala 122:34]
  wire [31:0] _out_bits_addr_T_5 = _out_bits_addr_T | _GEN_25; // @[Fragmenter.scala 122:34]
  wire  irr_valid = deq_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_2 = auto_out_arready & irr_valid; // @[Decoupled.scala 40:37]
  wire [8:0] _GEN_26 = {{1'd0}, len}; // @[Fragmenter.scala 127:25]
  wire [8:0] _rlen_T_1 = _GEN_26 - beats; // @[Fragmenter.scala 127:25]
  wire [8:0] _GEN_4 = _T_2 ? _rlen_T_1 : {{1'd0}, r_len}; // @[Fragmenter.scala 124:27 Fragmenter.scala 127:18 Fragmenter.scala 62:25]
  reg  busy_1; // @[Fragmenter.scala 60:29]
  reg [31:0] r_addr_1; // @[Fragmenter.scala 61:25]
  reg [7:0] r_len_1; // @[Fragmenter.scala 62:25]
  wire [7:0] irr_1_bits_len = deq_1_io_deq_bits_len; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire [7:0] len_1 = busy_1 ? r_len_1 : irr_1_bits_len; // @[Fragmenter.scala 64:23]
  wire [31:0] irr_1_bits_addr = deq_1_io_deq_bits_addr; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire [31:0] addr_1 = busy_1 ? r_addr_1 : irr_1_bits_addr; // @[Fragmenter.scala 65:23]
  wire [7:0] alignment_1 = addr_1[10:3]; // @[Fragmenter.scala 69:29]
  wire [7:0] _GEN_27 = {{1'd0}, len_1[7:1]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_8 = len_1 | _GEN_27; // @[package.scala 253:43]
  wire [7:0] _GEN_28 = {{2'd0}, _fillLow_T_8[7:2]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_10 = _fillLow_T_8 | _GEN_28; // @[package.scala 253:43]
  wire [7:0] _GEN_29 = {{4'd0}, _fillLow_T_10[7:4]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_12 = _fillLow_T_10 | _GEN_29; // @[package.scala 253:43]
  wire [6:0] fillLow_1 = _fillLow_T_12[7:1]; // @[Fragmenter.scala 85:37]
  wire [7:0] _wipeHigh_T_11 = ~len_1; // @[Fragmenter.scala 86:32]
  wire [8:0] _wipeHigh_T_12 = {_wipeHigh_T_11, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_14 = _wipeHigh_T_11 | _wipeHigh_T_12[7:0]; // @[package.scala 244:43]
  wire [9:0] _wipeHigh_T_15 = {_wipeHigh_T_14, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_17 = _wipeHigh_T_14 | _wipeHigh_T_15[7:0]; // @[package.scala 244:43]
  wire [11:0] _wipeHigh_T_18 = {_wipeHigh_T_17, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_20 = _wipeHigh_T_17 | _wipeHigh_T_18[7:0]; // @[package.scala 244:43]
  wire [7:0] wipeHigh_1 = ~_wipeHigh_T_20; // @[Fragmenter.scala 86:24]
  wire [7:0] _GEN_30 = {{1'd0}, fillLow_1}; // @[Fragmenter.scala 87:32]
  wire [7:0] remain1_1 = _GEN_30 | wipeHigh_1; // @[Fragmenter.scala 87:32]
  wire [8:0] _align1_T_10 = {alignment_1, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_12 = alignment_1 | _align1_T_10[7:0]; // @[package.scala 244:43]
  wire [9:0] _align1_T_13 = {_align1_T_12, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_15 = _align1_T_12 | _align1_T_13[7:0]; // @[package.scala 244:43]
  wire [11:0] _align1_T_16 = {_align1_T_15, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_18 = _align1_T_15 | _align1_T_16[7:0]; // @[package.scala 244:43]
  wire [7:0] align1_1 = ~_align1_T_18; // @[Fragmenter.scala 88:24]
  wire [7:0] _maxSupported1_T_1 = remain1_1 & align1_1; // @[Fragmenter.scala 89:37]
  wire [7:0] maxSupported1_1 = _maxSupported1_T_1 & 8'h7; // @[Fragmenter.scala 89:46]
  wire [1:0] irr_1_bits_burst = deq_1_io_deq_bits_burst; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  fixed_1 = irr_1_bits_burst == 2'h0; // @[Fragmenter.scala 92:34]
  wire [2:0] irr_1_bits_size = deq_1_io_deq_bits_size; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  narrow_1 = irr_1_bits_size != 3'h3; // @[Fragmenter.scala 93:34]
  wire  bad_1 = fixed_1 | narrow_1; // @[Fragmenter.scala 94:25]
  wire [7:0] beats_lo_1 = bad_1 ? 8'h0 : maxSupported1_1; // @[Fragmenter.scala 97:25]
  wire [8:0] _beats_T_4 = {beats_lo_1, 1'h0}; // @[package.scala 232:35]
  wire [8:0] _beats_T_5 = _beats_T_4 | 9'h1; // @[package.scala 232:40]
  wire [8:0] _beats_T_6 = {1'h0,beats_lo_1}; // @[Cat.scala 30:58]
  wire [8:0] _beats_T_7 = ~_beats_T_6; // @[package.scala 232:53]
  wire [8:0] w_beats = _beats_T_5 & _beats_T_7; // @[package.scala 232:51]
  wire [15:0] _GEN_31 = {{7'd0}, w_beats}; // @[Fragmenter.scala 100:38]
  wire [15:0] _inc_addr_T_2 = _GEN_31 << irr_1_bits_size; // @[Fragmenter.scala 100:38]
  wire [31:0] _GEN_32 = {{16'd0}, _inc_addr_T_2}; // @[Fragmenter.scala 100:29]
  wire [31:0] inc_addr_1 = addr_1 + _GEN_32; // @[Fragmenter.scala 100:29]
  wire [15:0] _wrapMask_T_2 = {irr_1_bits_len,8'hff}; // @[Cat.scala 30:58]
  wire [22:0] _GEN_33 = {{7'd0}, _wrapMask_T_2}; // @[Bundles.scala 31:21]
  wire [22:0] _wrapMask_T_3 = _GEN_33 << irr_1_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] wrapMask_1 = _wrapMask_T_3[22:8]; // @[Bundles.scala 31:30]
  wire [31:0] _GEN_34 = {{17'd0}, wrapMask_1}; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_5 = inc_addr_1 & _GEN_34; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_6 = ~irr_1_bits_addr; // @[Fragmenter.scala 104:49]
  wire [31:0] _mux_addr_T_7 = _mux_addr_T_6 | _GEN_34; // @[Fragmenter.scala 104:62]
  wire [31:0] _mux_addr_T_8 = ~_mux_addr_T_7; // @[Fragmenter.scala 104:47]
  wire [31:0] _mux_addr_T_9 = _mux_addr_T_5 | _mux_addr_T_8; // @[Fragmenter.scala 104:45]
  wire  aw_last = beats_lo_1 == len_1; // @[Fragmenter.scala 110:27]
  reg [8:0] w_counter; // @[Fragmenter.scala 164:30]
  wire  w_idle = w_counter == 9'h0; // @[Fragmenter.scala 165:30]
  reg  wbeats_latched; // @[Fragmenter.scala 150:35]
  wire  _in_awready_T = w_idle | wbeats_latched; // @[Fragmenter.scala 158:52]
  wire  in_awready = auto_out_awready & (w_idle | wbeats_latched); // @[Fragmenter.scala 158:35]
  wire [31:0] _out_bits_addr_T_7 = ~addr_1; // @[Fragmenter.scala 122:28]
  wire [9:0] _out_bits_addr_T_9 = 10'h7 << irr_1_bits_size; // @[package.scala 234:77]
  wire [2:0] _out_bits_addr_T_11 = ~_out_bits_addr_T_9[2:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_36 = {{29'd0}, _out_bits_addr_T_11}; // @[Fragmenter.scala 122:34]
  wire [31:0] _out_bits_addr_T_12 = _out_bits_addr_T_7 | _GEN_36; // @[Fragmenter.scala 122:34]
  wire  irr_1_valid = deq_1_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_5 = in_awready & irr_1_valid; // @[Decoupled.scala 40:37]
  wire [8:0] _GEN_37 = {{1'd0}, len_1}; // @[Fragmenter.scala 127:25]
  wire [8:0] _rlen_T_3 = _GEN_37 - w_beats; // @[Fragmenter.scala 127:25]
  wire [8:0] _GEN_9 = _T_5 ? _rlen_T_3 : {{1'd0}, r_len_1}; // @[Fragmenter.scala 124:27 Fragmenter.scala 127:18 Fragmenter.scala 62:25]
  wire  wbeats_valid = irr_1_valid & ~wbeats_latched; // @[Fragmenter.scala 159:35]
  wire  _GEN_10 = wbeats_valid & w_idle | wbeats_latched; // @[Fragmenter.scala 153:43 Fragmenter.scala 153:60 Fragmenter.scala 150:35]
  wire  bundleOut_0_awvalid = irr_1_valid & _in_awready_T; // @[Fragmenter.scala 157:35]
  wire  _T_7 = auto_out_awready & bundleOut_0_awvalid; // @[Decoupled.scala 40:37]
  wire [8:0] _wtodo_T = wbeats_valid ? w_beats : 9'h0; // @[Fragmenter.scala 166:35]
  wire [8:0] w_todo = w_idle ? _wtodo_T : w_counter; // @[Fragmenter.scala 166:23]
  wire  w_last = w_todo == 9'h1; // @[Fragmenter.scala 167:27]
  wire  in_wvalid = in_wdeq_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _bundleOut_0_wvalid_T_1 = ~w_idle | wbeats_valid; // @[Fragmenter.scala 173:51]
  wire  bundleOut_0_wvalid = in_wvalid & (~w_idle | wbeats_valid); // @[Fragmenter.scala 173:33]
  wire  _wcounter_T = auto_out_wready & bundleOut_0_wvalid; // @[Decoupled.scala 40:37]
  wire [8:0] _GEN_38 = {{8'd0}, _wcounter_T}; // @[Fragmenter.scala 168:27]
  wire [8:0] _wcounter_T_2 = w_todo - _GEN_38; // @[Fragmenter.scala 168:27]
  wire  in_wlast = in_wdeq_io_deq_bits_last; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  bundleOut_0_bready = auto_in_bready | ~auto_out_becho_real_last; // @[Fragmenter.scala 189:33]
  reg [1:0] error_0; // @[Fragmenter.scala 192:26]
  reg [1:0] error_1; // @[Fragmenter.scala 192:26]
  wire [1:0] _GEN_13 = auto_out_bid ? error_1 : error_0; // @[Fragmenter.scala 193:41 Fragmenter.scala 193:41]
  wire [1:0] _T_22 = 2'h1 << auto_out_bid; // @[OneHot.scala 65:12]
  wire  _T_26 = bundleOut_0_bready & auto_out_bvalid; // @[Decoupled.scala 40:37]
  wire [1:0] _error_0_T = error_0 | auto_out_bresp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_1_T = error_1 | auto_out_bresp; // @[Fragmenter.scala 195:70]
  Queue_13 deq ( // @[Decoupled.scala 296:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_id(deq_io_enq_bits_id),
    .io_enq_bits_addr(deq_io_enq_bits_addr),
    .io_enq_bits_len(deq_io_enq_bits_len),
    .io_enq_bits_size(deq_io_enq_bits_size),
    .io_enq_bits_burst(deq_io_enq_bits_burst),
    .io_enq_bits_echo_extra_id(deq_io_enq_bits_echo_extra_id),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_id(deq_io_deq_bits_id),
    .io_deq_bits_addr(deq_io_deq_bits_addr),
    .io_deq_bits_len(deq_io_deq_bits_len),
    .io_deq_bits_size(deq_io_deq_bits_size),
    .io_deq_bits_burst(deq_io_deq_bits_burst),
    .io_deq_bits_echo_extra_id(deq_io_deq_bits_echo_extra_id)
  );
  Queue_13 deq_1 ( // @[Decoupled.scala 296:21]
    .clock(deq_1_clock),
    .reset(deq_1_reset),
    .io_enq_ready(deq_1_io_enq_ready),
    .io_enq_valid(deq_1_io_enq_valid),
    .io_enq_bits_id(deq_1_io_enq_bits_id),
    .io_enq_bits_addr(deq_1_io_enq_bits_addr),
    .io_enq_bits_len(deq_1_io_enq_bits_len),
    .io_enq_bits_size(deq_1_io_enq_bits_size),
    .io_enq_bits_burst(deq_1_io_enq_bits_burst),
    .io_enq_bits_echo_extra_id(deq_1_io_enq_bits_echo_extra_id),
    .io_deq_ready(deq_1_io_deq_ready),
    .io_deq_valid(deq_1_io_deq_valid),
    .io_deq_bits_id(deq_1_io_deq_bits_id),
    .io_deq_bits_addr(deq_1_io_deq_bits_addr),
    .io_deq_bits_len(deq_1_io_deq_bits_len),
    .io_deq_bits_size(deq_1_io_deq_bits_size),
    .io_deq_bits_burst(deq_1_io_deq_bits_burst),
    .io_deq_bits_echo_extra_id(deq_1_io_deq_bits_echo_extra_id)
  );
  Queue_15 in_wdeq ( // @[Decoupled.scala 296:21]
    .clock(in_wdeq_clock),
    .reset(in_wdeq_reset),
    .io_enq_ready(in_wdeq_io_enq_ready),
    .io_enq_valid(in_wdeq_io_enq_valid),
    .io_enq_bits_data(in_wdeq_io_enq_bits_data),
    .io_enq_bits_strb(in_wdeq_io_enq_bits_strb),
    .io_enq_bits_last(in_wdeq_io_enq_bits_last),
    .io_deq_ready(in_wdeq_io_deq_ready),
    .io_deq_valid(in_wdeq_io_deq_valid),
    .io_deq_bits_data(in_wdeq_io_deq_bits_data),
    .io_deq_bits_strb(in_wdeq_io_deq_bits_strb),
    .io_deq_bits_last(in_wdeq_io_deq_bits_last)
  );
  assign auto_in_awready = deq_1_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign auto_in_wready = in_wdeq_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign auto_in_bvalid = auto_out_bvalid & auto_out_becho_real_last; // @[Fragmenter.scala 188:33]
  assign auto_in_bid = auto_out_bid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bresp = auto_out_bresp | _GEN_13; // @[Fragmenter.scala 193:41]
  assign auto_in_becho_extra_id = auto_out_becho_extra_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_arready = deq_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign auto_in_rvalid = auto_out_rvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rid = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rdata = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rresp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_recho_extra_id = auto_out_recho_extra_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rlast = auto_out_rlast & auto_out_recho_real_last; // @[Fragmenter.scala 183:41]
  assign auto_out_awvalid = irr_1_valid & _in_awready_T; // @[Fragmenter.scala 157:35]
  assign auto_out_awid = deq_1_io_deq_bits_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awaddr = ~_out_bits_addr_T_12; // @[Fragmenter.scala 122:26]
  assign auto_out_awlen = bad_1 ? 8'h0 : maxSupported1_1; // @[Fragmenter.scala 97:25]
  assign auto_out_awsize = deq_1_io_deq_bits_size; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awecho_extra_id = deq_1_io_deq_bits_echo_extra_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awecho_real_last = beats_lo_1 == len_1; // @[Fragmenter.scala 110:27]
  assign auto_out_wvalid = in_wvalid & (~w_idle | wbeats_valid); // @[Fragmenter.scala 173:33]
  assign auto_out_wdata = in_wdeq_io_deq_bits_data; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_wstrb = in_wdeq_io_deq_bits_strb; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_wlast = w_todo == 9'h1; // @[Fragmenter.scala 167:27]
  assign auto_out_bready = auto_in_bready | ~auto_out_becho_real_last; // @[Fragmenter.scala 189:33]
  assign auto_out_arvalid = deq_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  assign auto_out_arid = deq_io_deq_bits_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_araddr = ~_out_bits_addr_T_5; // @[Fragmenter.scala 122:26]
  assign auto_out_arlen = bad ? 8'h0 : maxSupported1; // @[Fragmenter.scala 97:25]
  assign auto_out_arsize = deq_io_deq_bits_size; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_arecho_extra_id = deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_arecho_real_last = beats_lo == len; // @[Fragmenter.scala 110:27]
  assign auto_out_rready = auto_in_rready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = auto_in_arvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_id = auto_in_arid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_addr = auto_in_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_len = auto_in_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_size = auto_in_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_burst = auto_in_arburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_echo_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_deq_ready = auto_out_arready & ar_last; // @[Fragmenter.scala 111:30]
  assign deq_1_clock = clock;
  assign deq_1_reset = reset;
  assign deq_1_io_enq_valid = auto_in_awvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_id = auto_in_awid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_addr = auto_in_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_len = auto_in_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_size = auto_in_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_burst = auto_in_awburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_echo_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_deq_ready = in_awready & aw_last; // @[Fragmenter.scala 111:30]
  assign in_wdeq_clock = clock;
  assign in_wdeq_reset = reset;
  assign in_wdeq_io_enq_valid = auto_in_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_wdeq_io_enq_bits_data = auto_in_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_wdeq_io_enq_bits_strb = auto_in_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_wdeq_io_enq_bits_last = auto_in_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_wdeq_io_deq_ready = auto_out_wready & _bundleOut_0_wvalid_T_1; // @[Fragmenter.scala 174:33]
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 60:29]
      busy <= 1'h0; // @[Fragmenter.scala 60:29]
    end else if (_T_2) begin // @[Fragmenter.scala 124:27]
      busy <= ~ar_last; // @[Fragmenter.scala 125:16]
    end
    if (_T_2) begin // @[Fragmenter.scala 124:27]
      if (fixed) begin // @[Fragmenter.scala 106:60]
        r_addr <= irr_bits_addr; // @[Fragmenter.scala 107:20]
      end else if (irr_bits_burst == 2'h2) begin // @[Fragmenter.scala 103:59]
        r_addr <= _mux_addr_T_4; // @[Fragmenter.scala 104:20]
      end else begin
        r_addr <= inc_addr;
      end
    end
    r_len <= _GEN_4[7:0];
    if (reset) begin // @[Fragmenter.scala 60:29]
      busy_1 <= 1'h0; // @[Fragmenter.scala 60:29]
    end else if (_T_5) begin // @[Fragmenter.scala 124:27]
      busy_1 <= ~aw_last; // @[Fragmenter.scala 125:16]
    end
    if (_T_5) begin // @[Fragmenter.scala 124:27]
      if (fixed_1) begin // @[Fragmenter.scala 106:60]
        r_addr_1 <= irr_1_bits_addr; // @[Fragmenter.scala 107:20]
      end else if (irr_1_bits_burst == 2'h2) begin // @[Fragmenter.scala 103:59]
        r_addr_1 <= _mux_addr_T_9; // @[Fragmenter.scala 104:20]
      end else begin
        r_addr_1 <= inc_addr_1;
      end
    end
    r_len_1 <= _GEN_9[7:0];
    if (reset) begin // @[Fragmenter.scala 164:30]
      w_counter <= 9'h0; // @[Fragmenter.scala 164:30]
    end else begin
      w_counter <= _wcounter_T_2; // @[Fragmenter.scala 168:17]
    end
    if (reset) begin // @[Fragmenter.scala 150:35]
      wbeats_latched <= 1'h0; // @[Fragmenter.scala 150:35]
    end else if (_T_7) begin // @[Fragmenter.scala 154:28]
      wbeats_latched <= 1'h0; // @[Fragmenter.scala 154:45]
    end else begin
      wbeats_latched <= _GEN_10;
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_0 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[0] & _T_26) begin // @[Fragmenter.scala 195:36]
      if (auto_out_becho_real_last) begin // @[Fragmenter.scala 195:48]
        error_0 <= 2'h0;
      end else begin
        error_0 <= _error_0_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_1 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[1] & _T_26) begin // @[Fragmenter.scala 195:36]
      if (auto_out_becho_real_last) begin // @[Fragmenter.scala 195:48]
        error_1 <= 2'h0;
      end else begin
        error_1 <= _error_1_T;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_wcounter_T | w_todo != 9'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:169 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n"
            ); // @[Fragmenter.scala 169:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_wcounter_T | w_todo != 9'h0 | reset)) begin
          $fatal; // @[Fragmenter.scala 169:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~bundleOut_0_wvalid | ~in_wlast | w_last | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:178 assert (!out.w.valid || !in_w.bits.last || w_last)\n"); // @[Fragmenter.scala 178:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~bundleOut_0_wvalid | ~in_wlast | w_last | reset)) begin
          $fatal; // @[Fragmenter.scala 178:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_len = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  busy_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_addr_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  r_len_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  w_counter = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  wbeats_latched = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  error_0 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  error_1 = _RAND_9[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4IdIndexer(
  output        auto_in_awready,
  input         auto_in_awvalid,
  input  [3:0]  auto_in_awid,
  input  [31:0] auto_in_awaddr,
  input  [7:0]  auto_in_awlen,
  input  [2:0]  auto_in_awsize,
  input  [1:0]  auto_in_awburst,
  output        auto_in_wready,
  input         auto_in_wvalid,
  input  [63:0] auto_in_wdata,
  input  [7:0]  auto_in_wstrb,
  input         auto_in_wlast,
  input         auto_in_bready,
  output        auto_in_bvalid,
  output [3:0]  auto_in_bid,
  output [1:0]  auto_in_bresp,
  output        auto_in_arready,
  input         auto_in_arvalid,
  input  [3:0]  auto_in_arid,
  input  [31:0] auto_in_araddr,
  input  [7:0]  auto_in_arlen,
  input  [2:0]  auto_in_arsize,
  input  [1:0]  auto_in_arburst,
  input         auto_in_rready,
  output        auto_in_rvalid,
  output [3:0]  auto_in_rid,
  output [63:0] auto_in_rdata,
  output [1:0]  auto_in_rresp,
  output        auto_in_rlast,
  input         auto_out_awready,
  output        auto_out_awvalid,
  output        auto_out_awid,
  output [31:0] auto_out_awaddr,
  output [7:0]  auto_out_awlen,
  output [2:0]  auto_out_awsize,
  output [1:0]  auto_out_awburst,
  output [2:0]  auto_out_awecho_extra_id,
  input         auto_out_wready,
  output        auto_out_wvalid,
  output [63:0] auto_out_wdata,
  output [7:0]  auto_out_wstrb,
  output        auto_out_wlast,
  output        auto_out_bready,
  input         auto_out_bvalid,
  input         auto_out_bid,
  input  [1:0]  auto_out_bresp,
  input  [2:0]  auto_out_becho_extra_id,
  input         auto_out_arready,
  output        auto_out_arvalid,
  output        auto_out_arid,
  output [31:0] auto_out_araddr,
  output [7:0]  auto_out_arlen,
  output [2:0]  auto_out_arsize,
  output [1:0]  auto_out_arburst,
  output [2:0]  auto_out_arecho_extra_id,
  output        auto_out_rready,
  input         auto_out_rvalid,
  input         auto_out_rid,
  input  [63:0] auto_out_rdata,
  input  [1:0]  auto_out_rresp,
  input  [2:0]  auto_out_recho_extra_id,
  input         auto_out_rlast
);
  assign auto_in_awready = auto_out_awready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_wready = auto_out_wready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bvalid = auto_out_bvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bid = {auto_out_becho_extra_id,auto_out_bid}; // @[Cat.scala 30:58]
  assign auto_in_bresp = auto_out_bresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_arready = auto_out_arready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rvalid = auto_out_rvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rid = {auto_out_recho_extra_id,auto_out_rid}; // @[Cat.scala 30:58]
  assign auto_in_rdata = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rresp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rlast = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_awvalid = auto_in_awvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awid = auto_in_awid[0]; // @[Nodes.scala 1207:84 BundleMap.scala 247:19]
  assign auto_out_awaddr = auto_in_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awlen = auto_in_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awsize = auto_in_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awburst = auto_in_awburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awecho_extra_id = auto_in_awid[3:1]; // @[IdIndexer.scala 71:56]
  assign auto_out_wvalid = auto_in_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wdata = auto_in_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wstrb = auto_in_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wlast = auto_in_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_bready = auto_in_bready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arvalid = auto_in_arvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arid = auto_in_arid[0]; // @[Nodes.scala 1207:84 BundleMap.scala 247:19]
  assign auto_out_araddr = auto_in_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arlen = auto_in_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arsize = auto_in_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arburst = auto_in_arburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arecho_extra_id = auto_in_arid[3:1]; // @[IdIndexer.scala 70:56]
  assign auto_out_rready = auto_in_rready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
endmodule
module QueueCompatibility_4(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [3:0] io_enq_bits_tl_state_size,
  input  [6:0] io_enq_bits_tl_state_source,
  input        io_enq_bits_extra_id,
  input        io_deq_ready,
  output       io_deq_valid,
  output [3:0] io_deq_bits_tl_state_size,
  output [6:0] io_deq_bits_tl_state_source,
  output       io_deq_bits_extra_id
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:16]; // @[Decoupled.scala 218:16]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [4:0] ram_tl_state_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire [4:0] ram_tl_state_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_tl_state_source [0:16]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [4:0] ram_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_tl_state_source_MPORT_data; // @[Decoupled.scala 218:16]
  wire [4:0] ram_tl_state_source_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_source_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_source_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_extra_id [0:16]; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [4:0] ram_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [4:0] ram_extra_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [4:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 5'h10; // @[Counter.scala 72:24]
  wire [4:0] _value_T_1 = enq_ptr_value + 5'h1; // @[Counter.scala 76:24]
  wire  wrap_1 = deq_ptr_value == 5'h10; // @[Counter.scala 72:24]
  wire [4:0] _value_T_3 = deq_ptr_value + 5'h1; // @[Counter.scala 76:24]
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size_io_deq_bits_MPORT_addr >= 5'h11 ? _RAND_1[3:0] :
    ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = enq_ptr_value;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source_io_deq_bits_MPORT_addr >= 5'h11 ? _RAND_3[6:0]
     : ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id_io_deq_bits_MPORT_addr >= 5'h11 ? _RAND_5[0:0] :
    ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_extra_id_MPORT_data = io_enq_bits_extra_id;
  assign ram_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_extra_id_MPORT_mask = 1'h1;
  assign ram_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_extra_id = ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_extra_id_MPORT_en & ram_extra_id_MPORT_mask) begin
      ram_extra_id[ram_extra_id_MPORT_addr] <= ram_extra_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 5'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      if (wrap) begin // @[Counter.scala 86:20]
        enq_ptr_value <= 5'h0; // @[Counter.scala 86:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 5'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      if (wrap_1) begin // @[Counter.scala 86:20]
        deq_ptr_value <= 5'h0; // @[Counter.scala 86:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    ram_extra_id[initvar] = _RAND_4[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enq_ptr_value = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  deq_ptr_value = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueCompatibility_11(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [3:0] io_enq_bits_tl_state_size,
  input  [6:0] io_enq_bits_tl_state_source,
  input        io_enq_bits_extra_id,
  input        io_deq_ready,
  output       io_deq_valid,
  output [3:0] io_deq_bits_tl_state_size,
  output [6:0] io_deq_bits_tl_state_source,
  output       io_deq_bits_extra_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[Decoupled.scala 218:16]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_tl_state_source [0:0]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_tl_state_source_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_source_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_source_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_tl_state_source_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_extra_id [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_extra_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_extra_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_extra_id_MPORT_data = io_enq_bits_extra_id;
  assign ram_extra_id_MPORT_addr = 1'h0;
  assign ram_extra_id_MPORT_mask = 1'h1;
  assign ram_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_extra_id = ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_extra_id_MPORT_en & ram_extra_id_MPORT_mask) begin
      ram_extra_id[ram_extra_id_MPORT_addr] <= ram_extra_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_extra_id[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4UserYanker_1(
  input         clock,
  input         reset,
  output        auto_in_awready,
  input         auto_in_awvalid,
  input  [3:0]  auto_in_awid,
  input  [31:0] auto_in_awaddr,
  input  [7:0]  auto_in_awlen,
  input  [2:0]  auto_in_awsize,
  input  [1:0]  auto_in_awburst,
  input  [3:0]  auto_in_awecho_tl_state_size,
  input  [6:0]  auto_in_awecho_tl_state_source,
  input         auto_in_awecho_extra_id,
  output        auto_in_wready,
  input         auto_in_wvalid,
  input  [63:0] auto_in_wdata,
  input  [7:0]  auto_in_wstrb,
  input         auto_in_wlast,
  input         auto_in_bready,
  output        auto_in_bvalid,
  output [3:0]  auto_in_bid,
  output [1:0]  auto_in_bresp,
  output [3:0]  auto_in_becho_tl_state_size,
  output [6:0]  auto_in_becho_tl_state_source,
  output        auto_in_becho_extra_id,
  output        auto_in_arready,
  input         auto_in_arvalid,
  input  [3:0]  auto_in_arid,
  input  [31:0] auto_in_araddr,
  input  [7:0]  auto_in_arlen,
  input  [2:0]  auto_in_arsize,
  input  [1:0]  auto_in_arburst,
  input  [3:0]  auto_in_arecho_tl_state_size,
  input  [6:0]  auto_in_arecho_tl_state_source,
  input         auto_in_arecho_extra_id,
  input         auto_in_rready,
  output        auto_in_rvalid,
  output [3:0]  auto_in_rid,
  output [63:0] auto_in_rdata,
  output [1:0]  auto_in_rresp,
  output [3:0]  auto_in_recho_tl_state_size,
  output [6:0]  auto_in_recho_tl_state_source,
  output        auto_in_recho_extra_id,
  output        auto_in_rlast,
  input         auto_out_awready,
  output        auto_out_awvalid,
  output [3:0]  auto_out_awid,
  output [31:0] auto_out_awaddr,
  output [7:0]  auto_out_awlen,
  output [2:0]  auto_out_awsize,
  output [1:0]  auto_out_awburst,
  input         auto_out_wready,
  output        auto_out_wvalid,
  output [63:0] auto_out_wdata,
  output [7:0]  auto_out_wstrb,
  output        auto_out_wlast,
  output        auto_out_bready,
  input         auto_out_bvalid,
  input  [3:0]  auto_out_bid,
  input  [1:0]  auto_out_bresp,
  input         auto_out_arready,
  output        auto_out_arvalid,
  output [3:0]  auto_out_arid,
  output [31:0] auto_out_araddr,
  output [7:0]  auto_out_arlen,
  output [2:0]  auto_out_arsize,
  output [1:0]  auto_out_arburst,
  output        auto_out_rready,
  input         auto_out_rvalid,
  input  [3:0]  auto_out_rid,
  input  [63:0] auto_out_rdata,
  input  [1:0]  auto_out_rresp,
  input         auto_out_rlast
);
  wire  QueueCompatibility_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_1_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_1_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_1_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_2_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_2_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_2_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_3_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_3_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_3_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_4_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_4_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_4_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_5_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_5_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_5_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_6_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_6_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_6_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_7_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_7_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_7_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_8_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_8_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_8_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_8_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_9_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_9_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_9_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_9_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_10_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_10_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_10_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_10_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_11_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_11_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_11_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_11_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_12_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_12_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_12_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_12_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_13_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_13_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_13_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_13_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_14_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_14_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_14_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_14_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_15_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_15_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_15_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_15_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_16_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_16_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_16_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_16_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_17_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_17_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_17_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_17_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_18_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_18_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_18_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_18_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_19_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_19_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_19_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_19_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_20_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_20_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_20_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_20_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_21_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_21_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_21_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_21_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_22_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_22_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_22_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_22_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_23_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_23_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_23_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_23_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_24_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_24_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_24_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_24_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_25_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_25_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_25_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_25_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_26_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_26_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_26_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_26_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_27_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_27_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_27_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_27_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_28_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_28_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_28_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_28_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_29_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_29_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_29_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_29_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_30_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_30_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_30_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_30_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_31_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_31_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_31_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_31_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  _arready_WIRE_0 = QueueCompatibility_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _arready_WIRE_1 = QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_1 = 4'h1 == auto_in_arid ? _arready_WIRE_1 : _arready_WIRE_0; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_2 = QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_2 = 4'h2 == auto_in_arid ? _arready_WIRE_2 : _GEN_1; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_3 = QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_3 = 4'h3 == auto_in_arid ? _arready_WIRE_3 : _GEN_2; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_4 = QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_4 = 4'h4 == auto_in_arid ? _arready_WIRE_4 : _GEN_3; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_5 = QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_5 = 4'h5 == auto_in_arid ? _arready_WIRE_5 : _GEN_4; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_6 = QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_6 = 4'h6 == auto_in_arid ? _arready_WIRE_6 : _GEN_5; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_7 = QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_7 = 4'h7 == auto_in_arid ? _arready_WIRE_7 : _GEN_6; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_8 = QueueCompatibility_8_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_8 = 4'h8 == auto_in_arid ? _arready_WIRE_8 : _GEN_7; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_9 = QueueCompatibility_9_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_9 = 4'h9 == auto_in_arid ? _arready_WIRE_9 : _GEN_8; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_10 = QueueCompatibility_10_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_10 = 4'ha == auto_in_arid ? _arready_WIRE_10 : _GEN_9; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_11 = QueueCompatibility_11_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_11 = 4'hb == auto_in_arid ? _arready_WIRE_11 : _GEN_10; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_12 = QueueCompatibility_12_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_12 = 4'hc == auto_in_arid ? _arready_WIRE_12 : _GEN_11; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_13 = QueueCompatibility_13_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_13 = 4'hd == auto_in_arid ? _arready_WIRE_13 : _GEN_12; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_14 = QueueCompatibility_14_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_14 = 4'he == auto_in_arid ? _arready_WIRE_14 : _GEN_13; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _arready_WIRE_15 = QueueCompatibility_15_io_enq_ready; // @[UserYanker.scala 55:25 UserYanker.scala 55:25]
  wire  _GEN_15 = 4'hf == auto_in_arid ? _arready_WIRE_15 : _GEN_14; // @[UserYanker.scala 56:36 UserYanker.scala 56:36]
  wire  _rvalid_WIRE_0 = QueueCompatibility_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _rvalid_WIRE_1 = QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_17 = 4'h1 == auto_out_rid ? _rvalid_WIRE_1 : _rvalid_WIRE_0; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_2 = QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_18 = 4'h2 == auto_out_rid ? _rvalid_WIRE_2 : _GEN_17; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_3 = QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_19 = 4'h3 == auto_out_rid ? _rvalid_WIRE_3 : _GEN_18; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_4 = QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_20 = 4'h4 == auto_out_rid ? _rvalid_WIRE_4 : _GEN_19; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_5 = QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_21 = 4'h5 == auto_out_rid ? _rvalid_WIRE_5 : _GEN_20; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_6 = QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_22 = 4'h6 == auto_out_rid ? _rvalid_WIRE_6 : _GEN_21; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_7 = QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_23 = 4'h7 == auto_out_rid ? _rvalid_WIRE_7 : _GEN_22; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_8 = QueueCompatibility_8_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_24 = 4'h8 == auto_out_rid ? _rvalid_WIRE_8 : _GEN_23; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_9 = QueueCompatibility_9_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_25 = 4'h9 == auto_out_rid ? _rvalid_WIRE_9 : _GEN_24; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_10 = QueueCompatibility_10_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_26 = 4'ha == auto_out_rid ? _rvalid_WIRE_10 : _GEN_25; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_11 = QueueCompatibility_11_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_27 = 4'hb == auto_out_rid ? _rvalid_WIRE_11 : _GEN_26; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_12 = QueueCompatibility_12_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_28 = 4'hc == auto_out_rid ? _rvalid_WIRE_12 : _GEN_27; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_13 = QueueCompatibility_13_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_29 = 4'hd == auto_out_rid ? _rvalid_WIRE_13 : _GEN_28; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_14 = QueueCompatibility_14_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_30 = 4'he == auto_out_rid ? _rvalid_WIRE_14 : _GEN_29; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rvalid_WIRE_15 = QueueCompatibility_15_io_deq_valid; // @[UserYanker.scala 61:24 UserYanker.scala 61:24]
  wire  _GEN_31 = 4'hf == auto_out_rid ? _rvalid_WIRE_15 : _GEN_30; // @[UserYanker.scala 63:28 UserYanker.scala 63:28]
  wire  _rWIRE_0_extra_id = QueueCompatibility_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _rWIRE_1_extra_id = QueueCompatibility_1_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_33 = 4'h1 == auto_out_rid ? _rWIRE_1_extra_id : _rWIRE_0_extra_id; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_2_extra_id = QueueCompatibility_2_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_34 = 4'h2 == auto_out_rid ? _rWIRE_2_extra_id : _GEN_33; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_3_extra_id = QueueCompatibility_3_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_35 = 4'h3 == auto_out_rid ? _rWIRE_3_extra_id : _GEN_34; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_4_extra_id = QueueCompatibility_4_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_36 = 4'h4 == auto_out_rid ? _rWIRE_4_extra_id : _GEN_35; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_5_extra_id = QueueCompatibility_5_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_37 = 4'h5 == auto_out_rid ? _rWIRE_5_extra_id : _GEN_36; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_6_extra_id = QueueCompatibility_6_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_38 = 4'h6 == auto_out_rid ? _rWIRE_6_extra_id : _GEN_37; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_7_extra_id = QueueCompatibility_7_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_39 = 4'h7 == auto_out_rid ? _rWIRE_7_extra_id : _GEN_38; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_8_extra_id = QueueCompatibility_8_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_40 = 4'h8 == auto_out_rid ? _rWIRE_8_extra_id : _GEN_39; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_9_extra_id = QueueCompatibility_9_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_41 = 4'h9 == auto_out_rid ? _rWIRE_9_extra_id : _GEN_40; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_10_extra_id = QueueCompatibility_10_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_42 = 4'ha == auto_out_rid ? _rWIRE_10_extra_id : _GEN_41; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_11_extra_id = QueueCompatibility_11_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_43 = 4'hb == auto_out_rid ? _rWIRE_11_extra_id : _GEN_42; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_12_extra_id = QueueCompatibility_12_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_44 = 4'hc == auto_out_rid ? _rWIRE_12_extra_id : _GEN_43; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_13_extra_id = QueueCompatibility_13_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_45 = 4'hd == auto_out_rid ? _rWIRE_13_extra_id : _GEN_44; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_14_extra_id = QueueCompatibility_14_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire  _GEN_46 = 4'he == auto_out_rid ? _rWIRE_14_extra_id : _GEN_45; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _rWIRE_15_extra_id = QueueCompatibility_15_io_deq_bits_extra_id; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _rWIRE_0_tl_state_source = QueueCompatibility_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _rWIRE_1_tl_state_source = QueueCompatibility_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_49 = 4'h1 == auto_out_rid ? _rWIRE_1_tl_state_source : _rWIRE_0_tl_state_source; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_2_tl_state_source = QueueCompatibility_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_50 = 4'h2 == auto_out_rid ? _rWIRE_2_tl_state_source : _GEN_49; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_3_tl_state_source = QueueCompatibility_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_51 = 4'h3 == auto_out_rid ? _rWIRE_3_tl_state_source : _GEN_50; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_4_tl_state_source = QueueCompatibility_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_52 = 4'h4 == auto_out_rid ? _rWIRE_4_tl_state_source : _GEN_51; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_5_tl_state_source = QueueCompatibility_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_53 = 4'h5 == auto_out_rid ? _rWIRE_5_tl_state_source : _GEN_52; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_6_tl_state_source = QueueCompatibility_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_54 = 4'h6 == auto_out_rid ? _rWIRE_6_tl_state_source : _GEN_53; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_7_tl_state_source = QueueCompatibility_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_55 = 4'h7 == auto_out_rid ? _rWIRE_7_tl_state_source : _GEN_54; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_8_tl_state_source = QueueCompatibility_8_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_56 = 4'h8 == auto_out_rid ? _rWIRE_8_tl_state_source : _GEN_55; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_9_tl_state_source = QueueCompatibility_9_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_57 = 4'h9 == auto_out_rid ? _rWIRE_9_tl_state_source : _GEN_56; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_10_tl_state_source = QueueCompatibility_10_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_58 = 4'ha == auto_out_rid ? _rWIRE_10_tl_state_source : _GEN_57; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_11_tl_state_source = QueueCompatibility_11_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_59 = 4'hb == auto_out_rid ? _rWIRE_11_tl_state_source : _GEN_58; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_12_tl_state_source = QueueCompatibility_12_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_60 = 4'hc == auto_out_rid ? _rWIRE_12_tl_state_source : _GEN_59; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_13_tl_state_source = QueueCompatibility_13_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_61 = 4'hd == auto_out_rid ? _rWIRE_13_tl_state_source : _GEN_60; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_14_tl_state_source = QueueCompatibility_14_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [6:0] _GEN_62 = 4'he == auto_out_rid ? _rWIRE_14_tl_state_source : _GEN_61; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _rWIRE_15_tl_state_source = QueueCompatibility_15_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _rWIRE_0_tl_state_size = QueueCompatibility_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _rWIRE_1_tl_state_size = QueueCompatibility_1_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_65 = 4'h1 == auto_out_rid ? _rWIRE_1_tl_state_size : _rWIRE_0_tl_state_size; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_2_tl_state_size = QueueCompatibility_2_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_66 = 4'h2 == auto_out_rid ? _rWIRE_2_tl_state_size : _GEN_65; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_3_tl_state_size = QueueCompatibility_3_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_67 = 4'h3 == auto_out_rid ? _rWIRE_3_tl_state_size : _GEN_66; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_4_tl_state_size = QueueCompatibility_4_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_68 = 4'h4 == auto_out_rid ? _rWIRE_4_tl_state_size : _GEN_67; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_5_tl_state_size = QueueCompatibility_5_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_69 = 4'h5 == auto_out_rid ? _rWIRE_5_tl_state_size : _GEN_68; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_6_tl_state_size = QueueCompatibility_6_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_70 = 4'h6 == auto_out_rid ? _rWIRE_6_tl_state_size : _GEN_69; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_7_tl_state_size = QueueCompatibility_7_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_71 = 4'h7 == auto_out_rid ? _rWIRE_7_tl_state_size : _GEN_70; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_8_tl_state_size = QueueCompatibility_8_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_72 = 4'h8 == auto_out_rid ? _rWIRE_8_tl_state_size : _GEN_71; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_9_tl_state_size = QueueCompatibility_9_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_73 = 4'h9 == auto_out_rid ? _rWIRE_9_tl_state_size : _GEN_72; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_10_tl_state_size = QueueCompatibility_10_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_74 = 4'ha == auto_out_rid ? _rWIRE_10_tl_state_size : _GEN_73; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_11_tl_state_size = QueueCompatibility_11_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_75 = 4'hb == auto_out_rid ? _rWIRE_11_tl_state_size : _GEN_74; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_12_tl_state_size = QueueCompatibility_12_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_76 = 4'hc == auto_out_rid ? _rWIRE_12_tl_state_size : _GEN_75; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_13_tl_state_size = QueueCompatibility_13_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_77 = 4'hd == auto_out_rid ? _rWIRE_13_tl_state_size : _GEN_76; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_14_tl_state_size = QueueCompatibility_14_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [3:0] _GEN_78 = 4'he == auto_out_rid ? _rWIRE_14_tl_state_size : _GEN_77; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _rWIRE_15_tl_state_size = QueueCompatibility_15_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:23 UserYanker.scala 62:23]
  wire [15:0] _arsel_T = 16'h1 << auto_in_arid; // @[OneHot.scala 65:12]
  wire  arsel_0 = _arsel_T[0]; // @[UserYanker.scala 67:55]
  wire  arsel_1 = _arsel_T[1]; // @[UserYanker.scala 67:55]
  wire  arsel_2 = _arsel_T[2]; // @[UserYanker.scala 67:55]
  wire  arsel_3 = _arsel_T[3]; // @[UserYanker.scala 67:55]
  wire  arsel_4 = _arsel_T[4]; // @[UserYanker.scala 67:55]
  wire  arsel_5 = _arsel_T[5]; // @[UserYanker.scala 67:55]
  wire  arsel_6 = _arsel_T[6]; // @[UserYanker.scala 67:55]
  wire  arsel_7 = _arsel_T[7]; // @[UserYanker.scala 67:55]
  wire  arsel_8 = _arsel_T[8]; // @[UserYanker.scala 67:55]
  wire  arsel_9 = _arsel_T[9]; // @[UserYanker.scala 67:55]
  wire  arsel_10 = _arsel_T[10]; // @[UserYanker.scala 67:55]
  wire  arsel_11 = _arsel_T[11]; // @[UserYanker.scala 67:55]
  wire  arsel_12 = _arsel_T[12]; // @[UserYanker.scala 67:55]
  wire  arsel_13 = _arsel_T[13]; // @[UserYanker.scala 67:55]
  wire  arsel_14 = _arsel_T[14]; // @[UserYanker.scala 67:55]
  wire  arsel_15 = _arsel_T[15]; // @[UserYanker.scala 67:55]
  wire [15:0] _rsel_T = 16'h1 << auto_out_rid; // @[OneHot.scala 65:12]
  wire  rsel_0 = _rsel_T[0]; // @[UserYanker.scala 68:55]
  wire  rsel_1 = _rsel_T[1]; // @[UserYanker.scala 68:55]
  wire  rsel_2 = _rsel_T[2]; // @[UserYanker.scala 68:55]
  wire  rsel_3 = _rsel_T[3]; // @[UserYanker.scala 68:55]
  wire  rsel_4 = _rsel_T[4]; // @[UserYanker.scala 68:55]
  wire  rsel_5 = _rsel_T[5]; // @[UserYanker.scala 68:55]
  wire  rsel_6 = _rsel_T[6]; // @[UserYanker.scala 68:55]
  wire  rsel_7 = _rsel_T[7]; // @[UserYanker.scala 68:55]
  wire  rsel_8 = _rsel_T[8]; // @[UserYanker.scala 68:55]
  wire  rsel_9 = _rsel_T[9]; // @[UserYanker.scala 68:55]
  wire  rsel_10 = _rsel_T[10]; // @[UserYanker.scala 68:55]
  wire  rsel_11 = _rsel_T[11]; // @[UserYanker.scala 68:55]
  wire  rsel_12 = _rsel_T[12]; // @[UserYanker.scala 68:55]
  wire  rsel_13 = _rsel_T[13]; // @[UserYanker.scala 68:55]
  wire  rsel_14 = _rsel_T[14]; // @[UserYanker.scala 68:55]
  wire  rsel_15 = _rsel_T[15]; // @[UserYanker.scala 68:55]
  wire  _awready_WIRE_0 = QueueCompatibility_16_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _awready_WIRE_1 = QueueCompatibility_17_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_81 = 4'h1 == auto_in_awid ? _awready_WIRE_1 : _awready_WIRE_0; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_2 = QueueCompatibility_18_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_82 = 4'h2 == auto_in_awid ? _awready_WIRE_2 : _GEN_81; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_3 = QueueCompatibility_19_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_83 = 4'h3 == auto_in_awid ? _awready_WIRE_3 : _GEN_82; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_4 = QueueCompatibility_20_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_84 = 4'h4 == auto_in_awid ? _awready_WIRE_4 : _GEN_83; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_5 = QueueCompatibility_21_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_85 = 4'h5 == auto_in_awid ? _awready_WIRE_5 : _GEN_84; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_6 = QueueCompatibility_22_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_86 = 4'h6 == auto_in_awid ? _awready_WIRE_6 : _GEN_85; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_7 = QueueCompatibility_23_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_87 = 4'h7 == auto_in_awid ? _awready_WIRE_7 : _GEN_86; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_8 = QueueCompatibility_24_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_88 = 4'h8 == auto_in_awid ? _awready_WIRE_8 : _GEN_87; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_9 = QueueCompatibility_25_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_89 = 4'h9 == auto_in_awid ? _awready_WIRE_9 : _GEN_88; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_10 = QueueCompatibility_26_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_90 = 4'ha == auto_in_awid ? _awready_WIRE_10 : _GEN_89; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_11 = QueueCompatibility_27_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_91 = 4'hb == auto_in_awid ? _awready_WIRE_11 : _GEN_90; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_12 = QueueCompatibility_28_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_92 = 4'hc == auto_in_awid ? _awready_WIRE_12 : _GEN_91; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_13 = QueueCompatibility_29_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_93 = 4'hd == auto_in_awid ? _awready_WIRE_13 : _GEN_92; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_14 = QueueCompatibility_30_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_94 = 4'he == auto_in_awid ? _awready_WIRE_14 : _GEN_93; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _awready_WIRE_15 = QueueCompatibility_31_io_enq_ready; // @[UserYanker.scala 76:25 UserYanker.scala 76:25]
  wire  _GEN_95 = 4'hf == auto_in_awid ? _awready_WIRE_15 : _GEN_94; // @[UserYanker.scala 77:36 UserYanker.scala 77:36]
  wire  _bvalid_WIRE_0 = QueueCompatibility_16_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _bvalid_WIRE_1 = QueueCompatibility_17_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_97 = 4'h1 == auto_out_bid ? _bvalid_WIRE_1 : _bvalid_WIRE_0; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_2 = QueueCompatibility_18_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_98 = 4'h2 == auto_out_bid ? _bvalid_WIRE_2 : _GEN_97; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_3 = QueueCompatibility_19_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_99 = 4'h3 == auto_out_bid ? _bvalid_WIRE_3 : _GEN_98; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_4 = QueueCompatibility_20_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_100 = 4'h4 == auto_out_bid ? _bvalid_WIRE_4 : _GEN_99; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_5 = QueueCompatibility_21_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_101 = 4'h5 == auto_out_bid ? _bvalid_WIRE_5 : _GEN_100; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_6 = QueueCompatibility_22_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_102 = 4'h6 == auto_out_bid ? _bvalid_WIRE_6 : _GEN_101; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_7 = QueueCompatibility_23_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_103 = 4'h7 == auto_out_bid ? _bvalid_WIRE_7 : _GEN_102; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_8 = QueueCompatibility_24_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_104 = 4'h8 == auto_out_bid ? _bvalid_WIRE_8 : _GEN_103; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_9 = QueueCompatibility_25_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_105 = 4'h9 == auto_out_bid ? _bvalid_WIRE_9 : _GEN_104; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_10 = QueueCompatibility_26_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_106 = 4'ha == auto_out_bid ? _bvalid_WIRE_10 : _GEN_105; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_11 = QueueCompatibility_27_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_107 = 4'hb == auto_out_bid ? _bvalid_WIRE_11 : _GEN_106; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_12 = QueueCompatibility_28_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_108 = 4'hc == auto_out_bid ? _bvalid_WIRE_12 : _GEN_107; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_13 = QueueCompatibility_29_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_109 = 4'hd == auto_out_bid ? _bvalid_WIRE_13 : _GEN_108; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_14 = QueueCompatibility_30_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_110 = 4'he == auto_out_bid ? _bvalid_WIRE_14 : _GEN_109; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bvalid_WIRE_15 = QueueCompatibility_31_io_deq_valid; // @[UserYanker.scala 82:24 UserYanker.scala 82:24]
  wire  _GEN_111 = 4'hf == auto_out_bid ? _bvalid_WIRE_15 : _GEN_110; // @[UserYanker.scala 84:28 UserYanker.scala 84:28]
  wire  _bWIRE_0_extra_id = QueueCompatibility_16_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _bWIRE_1_extra_id = QueueCompatibility_17_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_113 = 4'h1 == auto_out_bid ? _bWIRE_1_extra_id : _bWIRE_0_extra_id; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_2_extra_id = QueueCompatibility_18_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_114 = 4'h2 == auto_out_bid ? _bWIRE_2_extra_id : _GEN_113; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_3_extra_id = QueueCompatibility_19_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_115 = 4'h3 == auto_out_bid ? _bWIRE_3_extra_id : _GEN_114; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_4_extra_id = QueueCompatibility_20_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_116 = 4'h4 == auto_out_bid ? _bWIRE_4_extra_id : _GEN_115; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_5_extra_id = QueueCompatibility_21_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_117 = 4'h5 == auto_out_bid ? _bWIRE_5_extra_id : _GEN_116; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_6_extra_id = QueueCompatibility_22_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_118 = 4'h6 == auto_out_bid ? _bWIRE_6_extra_id : _GEN_117; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_7_extra_id = QueueCompatibility_23_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_119 = 4'h7 == auto_out_bid ? _bWIRE_7_extra_id : _GEN_118; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_8_extra_id = QueueCompatibility_24_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_120 = 4'h8 == auto_out_bid ? _bWIRE_8_extra_id : _GEN_119; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_9_extra_id = QueueCompatibility_25_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_121 = 4'h9 == auto_out_bid ? _bWIRE_9_extra_id : _GEN_120; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_10_extra_id = QueueCompatibility_26_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_122 = 4'ha == auto_out_bid ? _bWIRE_10_extra_id : _GEN_121; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_11_extra_id = QueueCompatibility_27_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_123 = 4'hb == auto_out_bid ? _bWIRE_11_extra_id : _GEN_122; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_12_extra_id = QueueCompatibility_28_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_124 = 4'hc == auto_out_bid ? _bWIRE_12_extra_id : _GEN_123; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_13_extra_id = QueueCompatibility_29_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_125 = 4'hd == auto_out_bid ? _bWIRE_13_extra_id : _GEN_124; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_14_extra_id = QueueCompatibility_30_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire  _GEN_126 = 4'he == auto_out_bid ? _bWIRE_14_extra_id : _GEN_125; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire  _bWIRE_15_extra_id = QueueCompatibility_31_io_deq_bits_extra_id; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _bWIRE_0_tl_state_source = QueueCompatibility_16_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _bWIRE_1_tl_state_source = QueueCompatibility_17_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_129 = 4'h1 == auto_out_bid ? _bWIRE_1_tl_state_source : _bWIRE_0_tl_state_source; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_2_tl_state_source = QueueCompatibility_18_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_130 = 4'h2 == auto_out_bid ? _bWIRE_2_tl_state_source : _GEN_129; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_3_tl_state_source = QueueCompatibility_19_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_131 = 4'h3 == auto_out_bid ? _bWIRE_3_tl_state_source : _GEN_130; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_4_tl_state_source = QueueCompatibility_20_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_132 = 4'h4 == auto_out_bid ? _bWIRE_4_tl_state_source : _GEN_131; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_5_tl_state_source = QueueCompatibility_21_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_133 = 4'h5 == auto_out_bid ? _bWIRE_5_tl_state_source : _GEN_132; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_6_tl_state_source = QueueCompatibility_22_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_134 = 4'h6 == auto_out_bid ? _bWIRE_6_tl_state_source : _GEN_133; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_7_tl_state_source = QueueCompatibility_23_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_135 = 4'h7 == auto_out_bid ? _bWIRE_7_tl_state_source : _GEN_134; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_8_tl_state_source = QueueCompatibility_24_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_136 = 4'h8 == auto_out_bid ? _bWIRE_8_tl_state_source : _GEN_135; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_9_tl_state_source = QueueCompatibility_25_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_137 = 4'h9 == auto_out_bid ? _bWIRE_9_tl_state_source : _GEN_136; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_10_tl_state_source = QueueCompatibility_26_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_138 = 4'ha == auto_out_bid ? _bWIRE_10_tl_state_source : _GEN_137; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_11_tl_state_source = QueueCompatibility_27_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_139 = 4'hb == auto_out_bid ? _bWIRE_11_tl_state_source : _GEN_138; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_12_tl_state_source = QueueCompatibility_28_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_140 = 4'hc == auto_out_bid ? _bWIRE_12_tl_state_source : _GEN_139; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_13_tl_state_source = QueueCompatibility_29_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_141 = 4'hd == auto_out_bid ? _bWIRE_13_tl_state_source : _GEN_140; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_14_tl_state_source = QueueCompatibility_30_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [6:0] _GEN_142 = 4'he == auto_out_bid ? _bWIRE_14_tl_state_source : _GEN_141; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [6:0] _bWIRE_15_tl_state_source = QueueCompatibility_31_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _bWIRE_0_tl_state_size = QueueCompatibility_16_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _bWIRE_1_tl_state_size = QueueCompatibility_17_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_145 = 4'h1 == auto_out_bid ? _bWIRE_1_tl_state_size : _bWIRE_0_tl_state_size; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_2_tl_state_size = QueueCompatibility_18_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_146 = 4'h2 == auto_out_bid ? _bWIRE_2_tl_state_size : _GEN_145; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_3_tl_state_size = QueueCompatibility_19_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_147 = 4'h3 == auto_out_bid ? _bWIRE_3_tl_state_size : _GEN_146; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_4_tl_state_size = QueueCompatibility_20_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_148 = 4'h4 == auto_out_bid ? _bWIRE_4_tl_state_size : _GEN_147; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_5_tl_state_size = QueueCompatibility_21_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_149 = 4'h5 == auto_out_bid ? _bWIRE_5_tl_state_size : _GEN_148; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_6_tl_state_size = QueueCompatibility_22_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_150 = 4'h6 == auto_out_bid ? _bWIRE_6_tl_state_size : _GEN_149; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_7_tl_state_size = QueueCompatibility_23_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_151 = 4'h7 == auto_out_bid ? _bWIRE_7_tl_state_size : _GEN_150; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_8_tl_state_size = QueueCompatibility_24_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_152 = 4'h8 == auto_out_bid ? _bWIRE_8_tl_state_size : _GEN_151; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_9_tl_state_size = QueueCompatibility_25_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_153 = 4'h9 == auto_out_bid ? _bWIRE_9_tl_state_size : _GEN_152; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_10_tl_state_size = QueueCompatibility_26_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_154 = 4'ha == auto_out_bid ? _bWIRE_10_tl_state_size : _GEN_153; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_11_tl_state_size = QueueCompatibility_27_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_155 = 4'hb == auto_out_bid ? _bWIRE_11_tl_state_size : _GEN_154; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_12_tl_state_size = QueueCompatibility_28_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_156 = 4'hc == auto_out_bid ? _bWIRE_12_tl_state_size : _GEN_155; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_13_tl_state_size = QueueCompatibility_29_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_157 = 4'hd == auto_out_bid ? _bWIRE_13_tl_state_size : _GEN_156; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_14_tl_state_size = QueueCompatibility_30_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [3:0] _GEN_158 = 4'he == auto_out_bid ? _bWIRE_14_tl_state_size : _GEN_157; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  wire [3:0] _bWIRE_15_tl_state_size = QueueCompatibility_31_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:23 UserYanker.scala 83:23]
  wire [15:0] _awsel_T = 16'h1 << auto_in_awid; // @[OneHot.scala 65:12]
  wire  awsel_0 = _awsel_T[0]; // @[UserYanker.scala 88:55]
  wire  awsel_1 = _awsel_T[1]; // @[UserYanker.scala 88:55]
  wire  awsel_2 = _awsel_T[2]; // @[UserYanker.scala 88:55]
  wire  awsel_3 = _awsel_T[3]; // @[UserYanker.scala 88:55]
  wire  awsel_4 = _awsel_T[4]; // @[UserYanker.scala 88:55]
  wire  awsel_5 = _awsel_T[5]; // @[UserYanker.scala 88:55]
  wire  awsel_6 = _awsel_T[6]; // @[UserYanker.scala 88:55]
  wire  awsel_7 = _awsel_T[7]; // @[UserYanker.scala 88:55]
  wire  awsel_8 = _awsel_T[8]; // @[UserYanker.scala 88:55]
  wire  awsel_9 = _awsel_T[9]; // @[UserYanker.scala 88:55]
  wire  awsel_10 = _awsel_T[10]; // @[UserYanker.scala 88:55]
  wire  awsel_11 = _awsel_T[11]; // @[UserYanker.scala 88:55]
  wire  awsel_12 = _awsel_T[12]; // @[UserYanker.scala 88:55]
  wire  awsel_13 = _awsel_T[13]; // @[UserYanker.scala 88:55]
  wire  awsel_14 = _awsel_T[14]; // @[UserYanker.scala 88:55]
  wire  awsel_15 = _awsel_T[15]; // @[UserYanker.scala 88:55]
  wire [15:0] _bsel_T = 16'h1 << auto_out_bid; // @[OneHot.scala 65:12]
  wire  bsel_0 = _bsel_T[0]; // @[UserYanker.scala 89:55]
  wire  bsel_1 = _bsel_T[1]; // @[UserYanker.scala 89:55]
  wire  bsel_2 = _bsel_T[2]; // @[UserYanker.scala 89:55]
  wire  bsel_3 = _bsel_T[3]; // @[UserYanker.scala 89:55]
  wire  bsel_4 = _bsel_T[4]; // @[UserYanker.scala 89:55]
  wire  bsel_5 = _bsel_T[5]; // @[UserYanker.scala 89:55]
  wire  bsel_6 = _bsel_T[6]; // @[UserYanker.scala 89:55]
  wire  bsel_7 = _bsel_T[7]; // @[UserYanker.scala 89:55]
  wire  bsel_8 = _bsel_T[8]; // @[UserYanker.scala 89:55]
  wire  bsel_9 = _bsel_T[9]; // @[UserYanker.scala 89:55]
  wire  bsel_10 = _bsel_T[10]; // @[UserYanker.scala 89:55]
  wire  bsel_11 = _bsel_T[11]; // @[UserYanker.scala 89:55]
  wire  bsel_12 = _bsel_T[12]; // @[UserYanker.scala 89:55]
  wire  bsel_13 = _bsel_T[13]; // @[UserYanker.scala 89:55]
  wire  bsel_14 = _bsel_T[14]; // @[UserYanker.scala 89:55]
  wire  bsel_15 = _bsel_T[15]; // @[UserYanker.scala 89:55]
  QueueCompatibility_4 QueueCompatibility ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_clock),
    .reset(QueueCompatibility_reset),
    .io_enq_ready(QueueCompatibility_io_enq_ready),
    .io_enq_valid(QueueCompatibility_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_io_deq_ready),
    .io_deq_valid(QueueCompatibility_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_1 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_1_clock),
    .reset(QueueCompatibility_1_reset),
    .io_enq_ready(QueueCompatibility_1_io_enq_ready),
    .io_enq_valid(QueueCompatibility_1_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_1_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_1_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_1_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_1_io_deq_ready),
    .io_deq_valid(QueueCompatibility_1_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_1_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_1_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_1_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_2 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_2_clock),
    .reset(QueueCompatibility_2_reset),
    .io_enq_ready(QueueCompatibility_2_io_enq_ready),
    .io_enq_valid(QueueCompatibility_2_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_2_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_2_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_2_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_2_io_deq_ready),
    .io_deq_valid(QueueCompatibility_2_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_2_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_2_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_2_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_3 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_3_clock),
    .reset(QueueCompatibility_3_reset),
    .io_enq_ready(QueueCompatibility_3_io_enq_ready),
    .io_enq_valid(QueueCompatibility_3_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_3_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_3_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_3_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_3_io_deq_ready),
    .io_deq_valid(QueueCompatibility_3_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_3_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_3_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_3_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_4 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_4_clock),
    .reset(QueueCompatibility_4_reset),
    .io_enq_ready(QueueCompatibility_4_io_enq_ready),
    .io_enq_valid(QueueCompatibility_4_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_4_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_4_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_4_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_4_io_deq_ready),
    .io_deq_valid(QueueCompatibility_4_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_4_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_4_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_4_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_5 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_5_clock),
    .reset(QueueCompatibility_5_reset),
    .io_enq_ready(QueueCompatibility_5_io_enq_ready),
    .io_enq_valid(QueueCompatibility_5_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_5_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_5_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_5_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_5_io_deq_ready),
    .io_deq_valid(QueueCompatibility_5_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_5_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_5_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_5_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_6 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_6_clock),
    .reset(QueueCompatibility_6_reset),
    .io_enq_ready(QueueCompatibility_6_io_enq_ready),
    .io_enq_valid(QueueCompatibility_6_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_6_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_6_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_6_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_6_io_deq_ready),
    .io_deq_valid(QueueCompatibility_6_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_6_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_6_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_6_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_7 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_7_clock),
    .reset(QueueCompatibility_7_reset),
    .io_enq_ready(QueueCompatibility_7_io_enq_ready),
    .io_enq_valid(QueueCompatibility_7_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_7_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_7_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_7_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_7_io_deq_ready),
    .io_deq_valid(QueueCompatibility_7_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_7_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_7_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_7_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_8 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_8_clock),
    .reset(QueueCompatibility_8_reset),
    .io_enq_ready(QueueCompatibility_8_io_enq_ready),
    .io_enq_valid(QueueCompatibility_8_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_8_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_8_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_8_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_8_io_deq_ready),
    .io_deq_valid(QueueCompatibility_8_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_8_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_8_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_8_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_9 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_9_clock),
    .reset(QueueCompatibility_9_reset),
    .io_enq_ready(QueueCompatibility_9_io_enq_ready),
    .io_enq_valid(QueueCompatibility_9_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_9_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_9_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_9_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_9_io_deq_ready),
    .io_deq_valid(QueueCompatibility_9_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_9_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_9_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_9_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_10 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_10_clock),
    .reset(QueueCompatibility_10_reset),
    .io_enq_ready(QueueCompatibility_10_io_enq_ready),
    .io_enq_valid(QueueCompatibility_10_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_10_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_10_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_10_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_10_io_deq_ready),
    .io_deq_valid(QueueCompatibility_10_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_10_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_10_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_10_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_11 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_11_clock),
    .reset(QueueCompatibility_11_reset),
    .io_enq_ready(QueueCompatibility_11_io_enq_ready),
    .io_enq_valid(QueueCompatibility_11_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_11_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_11_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_11_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_11_io_deq_ready),
    .io_deq_valid(QueueCompatibility_11_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_11_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_11_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_11_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_12 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_12_clock),
    .reset(QueueCompatibility_12_reset),
    .io_enq_ready(QueueCompatibility_12_io_enq_ready),
    .io_enq_valid(QueueCompatibility_12_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_12_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_12_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_12_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_12_io_deq_ready),
    .io_deq_valid(QueueCompatibility_12_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_12_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_12_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_12_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_13 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_13_clock),
    .reset(QueueCompatibility_13_reset),
    .io_enq_ready(QueueCompatibility_13_io_enq_ready),
    .io_enq_valid(QueueCompatibility_13_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_13_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_13_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_13_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_13_io_deq_ready),
    .io_deq_valid(QueueCompatibility_13_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_13_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_13_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_13_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_14 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_14_clock),
    .reset(QueueCompatibility_14_reset),
    .io_enq_ready(QueueCompatibility_14_io_enq_ready),
    .io_enq_valid(QueueCompatibility_14_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_14_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_14_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_14_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_14_io_deq_ready),
    .io_deq_valid(QueueCompatibility_14_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_14_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_14_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_14_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_15 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_15_clock),
    .reset(QueueCompatibility_15_reset),
    .io_enq_ready(QueueCompatibility_15_io_enq_ready),
    .io_enq_valid(QueueCompatibility_15_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_15_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_15_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_15_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_15_io_deq_ready),
    .io_deq_valid(QueueCompatibility_15_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_15_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_15_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_15_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_16 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_16_clock),
    .reset(QueueCompatibility_16_reset),
    .io_enq_ready(QueueCompatibility_16_io_enq_ready),
    .io_enq_valid(QueueCompatibility_16_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_16_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_16_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_16_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_16_io_deq_ready),
    .io_deq_valid(QueueCompatibility_16_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_16_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_16_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_16_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_17 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_17_clock),
    .reset(QueueCompatibility_17_reset),
    .io_enq_ready(QueueCompatibility_17_io_enq_ready),
    .io_enq_valid(QueueCompatibility_17_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_17_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_17_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_17_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_17_io_deq_ready),
    .io_deq_valid(QueueCompatibility_17_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_17_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_17_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_17_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_18 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_18_clock),
    .reset(QueueCompatibility_18_reset),
    .io_enq_ready(QueueCompatibility_18_io_enq_ready),
    .io_enq_valid(QueueCompatibility_18_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_18_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_18_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_18_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_18_io_deq_ready),
    .io_deq_valid(QueueCompatibility_18_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_18_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_18_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_18_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_19 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_19_clock),
    .reset(QueueCompatibility_19_reset),
    .io_enq_ready(QueueCompatibility_19_io_enq_ready),
    .io_enq_valid(QueueCompatibility_19_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_19_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_19_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_19_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_19_io_deq_ready),
    .io_deq_valid(QueueCompatibility_19_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_19_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_19_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_19_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_20 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_20_clock),
    .reset(QueueCompatibility_20_reset),
    .io_enq_ready(QueueCompatibility_20_io_enq_ready),
    .io_enq_valid(QueueCompatibility_20_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_20_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_20_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_20_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_20_io_deq_ready),
    .io_deq_valid(QueueCompatibility_20_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_20_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_20_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_20_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_21 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_21_clock),
    .reset(QueueCompatibility_21_reset),
    .io_enq_ready(QueueCompatibility_21_io_enq_ready),
    .io_enq_valid(QueueCompatibility_21_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_21_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_21_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_21_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_21_io_deq_ready),
    .io_deq_valid(QueueCompatibility_21_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_21_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_21_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_21_io_deq_bits_extra_id)
  );
  QueueCompatibility_4 QueueCompatibility_22 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_22_clock),
    .reset(QueueCompatibility_22_reset),
    .io_enq_ready(QueueCompatibility_22_io_enq_ready),
    .io_enq_valid(QueueCompatibility_22_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_22_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_22_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_22_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_22_io_deq_ready),
    .io_deq_valid(QueueCompatibility_22_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_22_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_22_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_22_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_23 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_23_clock),
    .reset(QueueCompatibility_23_reset),
    .io_enq_ready(QueueCompatibility_23_io_enq_ready),
    .io_enq_valid(QueueCompatibility_23_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_23_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_23_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_23_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_23_io_deq_ready),
    .io_deq_valid(QueueCompatibility_23_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_23_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_23_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_23_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_24 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_24_clock),
    .reset(QueueCompatibility_24_reset),
    .io_enq_ready(QueueCompatibility_24_io_enq_ready),
    .io_enq_valid(QueueCompatibility_24_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_24_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_24_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_24_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_24_io_deq_ready),
    .io_deq_valid(QueueCompatibility_24_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_24_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_24_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_24_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_25 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_25_clock),
    .reset(QueueCompatibility_25_reset),
    .io_enq_ready(QueueCompatibility_25_io_enq_ready),
    .io_enq_valid(QueueCompatibility_25_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_25_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_25_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_25_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_25_io_deq_ready),
    .io_deq_valid(QueueCompatibility_25_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_25_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_25_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_25_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_26 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_26_clock),
    .reset(QueueCompatibility_26_reset),
    .io_enq_ready(QueueCompatibility_26_io_enq_ready),
    .io_enq_valid(QueueCompatibility_26_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_26_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_26_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_26_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_26_io_deq_ready),
    .io_deq_valid(QueueCompatibility_26_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_26_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_26_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_26_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_27 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_27_clock),
    .reset(QueueCompatibility_27_reset),
    .io_enq_ready(QueueCompatibility_27_io_enq_ready),
    .io_enq_valid(QueueCompatibility_27_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_27_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_27_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_27_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_27_io_deq_ready),
    .io_deq_valid(QueueCompatibility_27_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_27_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_27_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_27_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_28 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_28_clock),
    .reset(QueueCompatibility_28_reset),
    .io_enq_ready(QueueCompatibility_28_io_enq_ready),
    .io_enq_valid(QueueCompatibility_28_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_28_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_28_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_28_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_28_io_deq_ready),
    .io_deq_valid(QueueCompatibility_28_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_28_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_28_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_28_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_29 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_29_clock),
    .reset(QueueCompatibility_29_reset),
    .io_enq_ready(QueueCompatibility_29_io_enq_ready),
    .io_enq_valid(QueueCompatibility_29_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_29_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_29_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_29_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_29_io_deq_ready),
    .io_deq_valid(QueueCompatibility_29_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_29_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_29_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_29_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_30 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_30_clock),
    .reset(QueueCompatibility_30_reset),
    .io_enq_ready(QueueCompatibility_30_io_enq_ready),
    .io_enq_valid(QueueCompatibility_30_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_30_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_30_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_30_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_30_io_deq_ready),
    .io_deq_valid(QueueCompatibility_30_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_30_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_30_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_30_io_deq_bits_extra_id)
  );
  QueueCompatibility_11 QueueCompatibility_31 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_31_clock),
    .reset(QueueCompatibility_31_reset),
    .io_enq_ready(QueueCompatibility_31_io_enq_ready),
    .io_enq_valid(QueueCompatibility_31_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_31_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_31_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_31_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_31_io_deq_ready),
    .io_deq_valid(QueueCompatibility_31_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_31_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_31_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_31_io_deq_bits_extra_id)
  );
  assign auto_in_awready = auto_out_awready & _GEN_95; // @[UserYanker.scala 77:36]
  assign auto_in_wready = auto_out_wready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bvalid = auto_out_bvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bid = auto_out_bid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bresp = auto_out_bresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_becho_tl_state_size = 4'hf == auto_out_bid ? _bWIRE_15_tl_state_size : _GEN_158; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_becho_tl_state_source = 4'hf == auto_out_bid ? _bWIRE_15_tl_state_source : _GEN_142; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_becho_extra_id = 4'hf == auto_out_bid ? _bWIRE_15_extra_id : _GEN_126; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_arready = auto_out_arready & _GEN_15; // @[UserYanker.scala 56:36]
  assign auto_in_rvalid = auto_out_rvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rid = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rdata = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rresp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_recho_tl_state_size = 4'hf == auto_out_rid ? _rWIRE_15_tl_state_size : _GEN_78; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_recho_tl_state_source = 4'hf == auto_out_rid ? _rWIRE_15_tl_state_source : _GEN_62; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_recho_extra_id = 4'hf == auto_out_rid ? _rWIRE_15_extra_id : _GEN_46; // @[BundleMap.scala 247:19 BundleMap.scala 247:19]
  assign auto_in_rlast = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_awvalid = auto_in_awvalid & _GEN_95; // @[UserYanker.scala 78:36]
  assign auto_out_awid = auto_in_awid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awaddr = auto_in_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awlen = auto_in_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awsize = auto_in_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awburst = auto_in_awburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wvalid = auto_in_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wdata = auto_in_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wstrb = auto_in_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wlast = auto_in_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_bready = auto_in_bready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arvalid = auto_in_arvalid & _GEN_15; // @[UserYanker.scala 57:36]
  assign auto_out_arid = auto_in_arid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_araddr = auto_in_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arlen = auto_in_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arsize = auto_in_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arburst = auto_in_arburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_rready = auto_in_rready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_clock = clock;
  assign QueueCompatibility_reset = reset;
  assign QueueCompatibility_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_0; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_0 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_1_clock = clock;
  assign QueueCompatibility_1_reset = reset;
  assign QueueCompatibility_1_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_1; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_1_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_1 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_2_clock = clock;
  assign QueueCompatibility_2_reset = reset;
  assign QueueCompatibility_2_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_2; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_2_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_2 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_3_clock = clock;
  assign QueueCompatibility_3_reset = reset;
  assign QueueCompatibility_3_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_3; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_3_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_3 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_4_clock = clock;
  assign QueueCompatibility_4_reset = reset;
  assign QueueCompatibility_4_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_4; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_4_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_4_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_4_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_4_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_4 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_5_clock = clock;
  assign QueueCompatibility_5_reset = reset;
  assign QueueCompatibility_5_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_5; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_5_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_5_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_5_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_5_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_5 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_6_clock = clock;
  assign QueueCompatibility_6_reset = reset;
  assign QueueCompatibility_6_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_6; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_6_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_6_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_6_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_6_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_6 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_7_clock = clock;
  assign QueueCompatibility_7_reset = reset;
  assign QueueCompatibility_7_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_7; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_7_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_7_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_7_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_7_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_7 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_8_clock = clock;
  assign QueueCompatibility_8_reset = reset;
  assign QueueCompatibility_8_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_8; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_8_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_8_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_8_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_8_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_8 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_9_clock = clock;
  assign QueueCompatibility_9_reset = reset;
  assign QueueCompatibility_9_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_9; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_9_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_9_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_9_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_9_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_9 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_10_clock = clock;
  assign QueueCompatibility_10_reset = reset;
  assign QueueCompatibility_10_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_10; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_10_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_10_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_10_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_10_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_10 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_11_clock = clock;
  assign QueueCompatibility_11_reset = reset;
  assign QueueCompatibility_11_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_11; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_11_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_11_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_11_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_11_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_11 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_12_clock = clock;
  assign QueueCompatibility_12_reset = reset;
  assign QueueCompatibility_12_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_12; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_12_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_12_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_12_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_12_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_12 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_13_clock = clock;
  assign QueueCompatibility_13_reset = reset;
  assign QueueCompatibility_13_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_13; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_13_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_13_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_13_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_13_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_13 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_14_clock = clock;
  assign QueueCompatibility_14_reset = reset;
  assign QueueCompatibility_14_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_14; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_14_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_14_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_14_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_14_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_14 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_15_clock = clock;
  assign QueueCompatibility_15_reset = reset;
  assign QueueCompatibility_15_io_enq_valid = auto_in_arvalid & auto_out_arready & arsel_15; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_15_io_enq_bits_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_15_io_enq_bits_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_15_io_enq_bits_extra_id = auto_in_arecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_15_io_deq_ready = auto_out_rvalid & auto_in_rready & rsel_15 & auto_out_rlast; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_16_clock = clock;
  assign QueueCompatibility_16_reset = reset;
  assign QueueCompatibility_16_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_0; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_16_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_16_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_16_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_16_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_0; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_17_clock = clock;
  assign QueueCompatibility_17_reset = reset;
  assign QueueCompatibility_17_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_1; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_17_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_17_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_17_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_17_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_1; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_18_clock = clock;
  assign QueueCompatibility_18_reset = reset;
  assign QueueCompatibility_18_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_2; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_18_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_18_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_18_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_18_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_2; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_19_clock = clock;
  assign QueueCompatibility_19_reset = reset;
  assign QueueCompatibility_19_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_3; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_19_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_19_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_19_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_19_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_3; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_20_clock = clock;
  assign QueueCompatibility_20_reset = reset;
  assign QueueCompatibility_20_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_4; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_20_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_20_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_20_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_20_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_4; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_21_clock = clock;
  assign QueueCompatibility_21_reset = reset;
  assign QueueCompatibility_21_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_5; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_21_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_21_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_21_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_21_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_5; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_22_clock = clock;
  assign QueueCompatibility_22_reset = reset;
  assign QueueCompatibility_22_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_6; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_22_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_22_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_22_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_22_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_6; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_23_clock = clock;
  assign QueueCompatibility_23_reset = reset;
  assign QueueCompatibility_23_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_7; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_23_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_23_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_23_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_23_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_7; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_24_clock = clock;
  assign QueueCompatibility_24_reset = reset;
  assign QueueCompatibility_24_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_8; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_24_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_24_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_24_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_24_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_8; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_25_clock = clock;
  assign QueueCompatibility_25_reset = reset;
  assign QueueCompatibility_25_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_9; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_25_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_25_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_25_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_25_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_9; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_26_clock = clock;
  assign QueueCompatibility_26_reset = reset;
  assign QueueCompatibility_26_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_10; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_26_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_26_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_26_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_26_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_10; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_27_clock = clock;
  assign QueueCompatibility_27_reset = reset;
  assign QueueCompatibility_27_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_11; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_27_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_27_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_27_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_27_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_11; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_28_clock = clock;
  assign QueueCompatibility_28_reset = reset;
  assign QueueCompatibility_28_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_12; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_28_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_28_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_28_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_28_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_12; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_29_clock = clock;
  assign QueueCompatibility_29_reset = reset;
  assign QueueCompatibility_29_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_13; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_29_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_29_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_29_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_29_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_13; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_30_clock = clock;
  assign QueueCompatibility_30_reset = reset;
  assign QueueCompatibility_30_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_14; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_30_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_30_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_30_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_30_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_14; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_31_clock = clock;
  assign QueueCompatibility_31_reset = reset;
  assign QueueCompatibility_31_io_enq_valid = auto_in_awvalid & auto_out_awready & awsel_15; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_31_io_enq_bits_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_31_io_enq_bits_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_31_io_enq_bits_extra_id = auto_in_awecho_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_31_io_deq_ready = auto_out_bvalid & auto_in_bready & bsel_15; // @[UserYanker.scala 91:53]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~auto_out_rvalid | _GEN_31 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:63 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 63:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_rvalid | _GEN_31 | reset)) begin
          $fatal; // @[UserYanker.scala 63:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~auto_out_bvalid | _GEN_111 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:84 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 84:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_bvalid | _GEN_111 | reset)) begin
          $fatal; // @[UserYanker.scala 84:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer_1(
  output        auto_in_awready,
  input         auto_in_awvalid,
  input  [4:0]  auto_in_awid,
  input  [31:0] auto_in_awaddr,
  input  [7:0]  auto_in_awlen,
  input  [2:0]  auto_in_awsize,
  input  [1:0]  auto_in_awburst,
  input  [3:0]  auto_in_awecho_tl_state_size,
  input  [6:0]  auto_in_awecho_tl_state_source,
  output        auto_in_wready,
  input         auto_in_wvalid,
  input  [63:0] auto_in_wdata,
  input  [7:0]  auto_in_wstrb,
  input         auto_in_wlast,
  input         auto_in_bready,
  output        auto_in_bvalid,
  output [4:0]  auto_in_bid,
  output [1:0]  auto_in_bresp,
  output [3:0]  auto_in_becho_tl_state_size,
  output [6:0]  auto_in_becho_tl_state_source,
  output        auto_in_arready,
  input         auto_in_arvalid,
  input  [4:0]  auto_in_arid,
  input  [31:0] auto_in_araddr,
  input  [7:0]  auto_in_arlen,
  input  [2:0]  auto_in_arsize,
  input  [1:0]  auto_in_arburst,
  input  [3:0]  auto_in_arecho_tl_state_size,
  input  [6:0]  auto_in_arecho_tl_state_source,
  input         auto_in_rready,
  output        auto_in_rvalid,
  output [4:0]  auto_in_rid,
  output [63:0] auto_in_rdata,
  output [1:0]  auto_in_rresp,
  output [3:0]  auto_in_recho_tl_state_size,
  output [6:0]  auto_in_recho_tl_state_source,
  output        auto_in_rlast,
  input         auto_out_awready,
  output        auto_out_awvalid,
  output [3:0]  auto_out_awid,
  output [31:0] auto_out_awaddr,
  output [7:0]  auto_out_awlen,
  output [2:0]  auto_out_awsize,
  output [1:0]  auto_out_awburst,
  output [3:0]  auto_out_awecho_tl_state_size,
  output [6:0]  auto_out_awecho_tl_state_source,
  output        auto_out_awecho_extra_id,
  input         auto_out_wready,
  output        auto_out_wvalid,
  output [63:0] auto_out_wdata,
  output [7:0]  auto_out_wstrb,
  output        auto_out_wlast,
  output        auto_out_bready,
  input         auto_out_bvalid,
  input  [3:0]  auto_out_bid,
  input  [1:0]  auto_out_bresp,
  input  [3:0]  auto_out_becho_tl_state_size,
  input  [6:0]  auto_out_becho_tl_state_source,
  input         auto_out_becho_extra_id,
  input         auto_out_arready,
  output        auto_out_arvalid,
  output [3:0]  auto_out_arid,
  output [31:0] auto_out_araddr,
  output [7:0]  auto_out_arlen,
  output [2:0]  auto_out_arsize,
  output [1:0]  auto_out_arburst,
  output [3:0]  auto_out_arecho_tl_state_size,
  output [6:0]  auto_out_arecho_tl_state_source,
  output        auto_out_arecho_extra_id,
  output        auto_out_rready,
  input         auto_out_rvalid,
  input  [3:0]  auto_out_rid,
  input  [63:0] auto_out_rdata,
  input  [1:0]  auto_out_rresp,
  input  [3:0]  auto_out_recho_tl_state_size,
  input  [6:0]  auto_out_recho_tl_state_source,
  input         auto_out_recho_extra_id,
  input         auto_out_rlast
);
  assign auto_in_awready = auto_out_awready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_wready = auto_out_wready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bvalid = auto_out_bvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bid = {auto_out_becho_extra_id,auto_out_bid}; // @[Cat.scala 30:58]
  assign auto_in_bresp = auto_out_bresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_becho_tl_state_size = auto_out_becho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_becho_tl_state_source = auto_out_becho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_arready = auto_out_arready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rvalid = auto_out_rvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rid = {auto_out_recho_extra_id,auto_out_rid}; // @[Cat.scala 30:58]
  assign auto_in_rdata = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rresp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_recho_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_recho_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rlast = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_awvalid = auto_in_awvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awid = auto_in_awid[3:0]; // @[Nodes.scala 1207:84 BundleMap.scala 247:19]
  assign auto_out_awaddr = auto_in_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awlen = auto_in_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awsize = auto_in_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awburst = auto_in_awburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awecho_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awecho_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awecho_extra_id = auto_in_awid[4]; // @[IdIndexer.scala 71:56]
  assign auto_out_wvalid = auto_in_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wdata = auto_in_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wstrb = auto_in_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wlast = auto_in_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_bready = auto_in_bready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arvalid = auto_in_arvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arid = auto_in_arid[3:0]; // @[Nodes.scala 1207:84 BundleMap.scala 247:19]
  assign auto_out_araddr = auto_in_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arlen = auto_in_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arsize = auto_in_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arburst = auto_in_arburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arecho_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arecho_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arecho_extra_id = auto_in_arid[4]; // @[IdIndexer.scala 70:56]
  assign auto_out_rready = auto_in_rready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
endmodule
module TLMonitor_10(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_a_bits_corrupt,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [2:0]  io_in_d_bits_size,
  input  [6:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [511:0] _RAND_12;
  reg [511:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [511:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_2 = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_3 = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_4 = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_5 = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_lo = mask_acc_2 | mask_size_2 & mask_eq_6; // @[Misc.scala 214:29]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_hi = mask_acc_2 | mask_size_2 & mask_eq_7; // @[Misc.scala 214:29]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_lo = mask_acc_3 | mask_size_2 & mask_eq_8; // @[Misc.scala 214:29]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_hi = mask_acc_3 | mask_size_2 & mask_eq_9; // @[Misc.scala 214:29]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_lo = mask_acc_4 | mask_size_2 & mask_eq_10; // @[Misc.scala 214:29]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_hi = mask_acc_4 | mask_size_2 & mask_eq_11; // @[Misc.scala 214:29]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_lo = mask_acc_5 | mask_size_2 & mask_eq_12; // @[Misc.scala 214:29]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_hi = mask_acc_5 | mask_size_2 & mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire [31:0] _T_180 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_181 = {1'b0,$signed(_T_180)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_183 = $signed(_T_181) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_184 = $signed(_T_183) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_185 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_186 = {1'b0,$signed(_T_185)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_188 = $signed(_T_186) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_189 = $signed(_T_188) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_190 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_191 = {1'b0,$signed(_T_190)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_193 = $signed(_T_191) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_194 = $signed(_T_193) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_195 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_196 = {1'b0,$signed(_T_195)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_198 = $signed(_T_196) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_199 = $signed(_T_198) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_200 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_201 = {1'b0,$signed(_T_200)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_203 = $signed(_T_201) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_204 = $signed(_T_203) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_208 = _T_184 | _T_189 | _T_194 | _T_199 | _T_204; // @[Parameters.scala 671:42]
  wire  _T_214 = ~reset; // @[Monitor.scala 42:11]
  wire  _T_264 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_266 = _source_ok_T_1 & _T_264; // @[Mux.scala 27:72]
  wire  _T_316 = _T_266 & _T_208; // @[Monitor.scala 83:78]
  wire  _T_330 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [7:0] _T_334 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_335 = _T_334 == 8'h0; // @[Monitor.scala 88:31]
  wire  _T_339 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18]
  wire  _T_343 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_559 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_572 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_669 = _T_264 & _T_208; // @[Parameters.scala 670:56]
  wire  _T_680 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_684 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_692 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_788 = source_ok & _T_669; // @[Monitor.scala 115:71]
  wire  _T_806 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [7:0] _T_916 = ~mask; // @[Monitor.scala 127:33]
  wire [7:0] _T_917 = io_in_a_bits_mask & _T_916; // @[Monitor.scala 127:31]
  wire  _T_918 = _T_917 == 8'h0; // @[Monitor.scala 127:40]
  wire  _T_922 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_1025 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_1033 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_1136 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_1144 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1247 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1259 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1263 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1267 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27]
  wire  _T_1275 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1279 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1283 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1311 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1331 = _T_1279 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1340 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1357 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1375 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [6:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_1405 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_1406 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_1410 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_1414 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_1418 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_1422 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [6:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_1429 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_1430 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_1438 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_1442 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_1450 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  reg [127:0] inflight; // @[Monitor.scala 611:27]
  reg [511:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [511:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  wire [8:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [9:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69]
  wire [511:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [511:0] _GEN_73 = {{496'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[511:1]}; // @[Monitor.scala 634:152]
  wire [511:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [511:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91]
  wire [511:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[511:1]}; // @[Monitor.scala 638:144]
  wire  _T_1456 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [127:0] _a_set_wo_ready_T = 128'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_1459 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [8:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [9:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [1026:0] _GEN_79 = {{1023'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [1026:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [1026:0] _GEN_81 = {{1023'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [1026:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [127:0] _T_1461 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_1463 = ~_T_1461[0]; // @[Monitor.scala 658:17]
  wire [127:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [1026:0] _GEN_19 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [1026:0] _GEN_20 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_1467 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_1469 = ~_T_1263; // @[Monitor.scala 671:74]
  wire  _T_1470 = io_in_d_valid & d_first_1 & ~_T_1263; // @[Monitor.scala 671:71]
  wire [127:0] _d_clr_wo_ready_T = 128'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1263 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [1038:0] _GEN_83 = {{1023'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [1038:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [127:0] d_clr = _d_first_T & d_first_1 & _T_1469 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [1038:0] _GEN_23 = _d_first_T & d_first_1 & _T_1469 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_1456 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [127:0] _T_1480 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_1482 = _T_1480[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_1487 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39]
  wire  _T_1488 = io_in_d_bits_opcode == _GEN_32 | _T_1487; // @[Monitor.scala 685:77]
  wire  _T_1492 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_1499 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_1500 = io_in_d_bits_opcode == _GEN_48 | _T_1499; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_1504 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_1514 = _T_1467 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_1469; // @[Monitor.scala 694:116]
  wire  _T_1516 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_1523 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [127:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [127:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [127:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [511:0] a_opcodes_set = _GEN_19[511:0];
  wire [511:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [511:0] d_opcodes_clr = _GEN_23[511:0];
  wire [511:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [511:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [511:0] a_sizes_set = _GEN_20[511:0];
  wire [511:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [511:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_1532 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [127:0] inflight_1; // @[Monitor.scala 723:35]
  reg [511:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25]
  wire [511:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [511:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93]
  wire [511:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[511:1]}; // @[Monitor.scala 747:146]
  wire  _T_1558 = io_in_d_valid & d_first_2 & _T_1263; // @[Monitor.scala 779:71]
  wire [127:0] d_clr_1 = _d_first_T & d_first_2 & _T_1263 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [1038:0] _GEN_68 = _d_first_T & d_first_2 & _T_1263 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire [127:0] _T_1566 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_1576 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36]
  wire [127:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [127:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [511:0] d_opcodes_clr_1 = _GEN_68[511:0];
  wire [511:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [511:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_1601 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 128'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 512'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 512'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 128'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 512'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_316 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_316 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_330 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_330 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_335 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_335 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_339 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_339 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_316 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_316 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_330 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_330 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_559 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_559 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_335 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_335 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_339 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_343 & ~(_T_339 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(_T_669 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(_T_669 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(_T_680 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(_T_680 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(_T_684 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(_T_684 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(_T_339 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_572 & ~(_T_339 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(_T_788 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(_T_788 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(_T_680 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(_T_680 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(_T_684 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_692 & ~(_T_684 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(_T_788 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(_T_788 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(_T_680 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(_T_680 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(_T_918 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_806 & ~(_T_918 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~(_T_1025 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~(_T_1025 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~(_T_684 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_922 & ~(_T_684 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~(_T_1136 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~(_T_1136 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~(_T_684 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1033 & ~(_T_684 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(_T_1247 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(_T_1247 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(_T_684 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(_T_684 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(_T_339 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1144 & ~(_T_339 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1259 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1259 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1263 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1263 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1263 & ~(_T_1267 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1263 & ~(_T_1267 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1263 & ~(_T_1275 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1263 & ~(_T_1275 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1263 & ~(_T_1279 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1263 & ~(_T_1279 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1283 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1283 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1283 & _T_214) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1283 & _T_214) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1283 & ~(_T_1267 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1283 & ~(_T_1267 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1283 & ~(_T_1275 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1283 & ~(_T_1275 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1311 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1311 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1311 & _T_214) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1311 & _T_214) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1311 & ~(_T_1267 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1311 & ~(_T_1267 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1311 & ~(_T_1331 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1311 & ~(_T_1331 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1340 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1340 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1340 & ~(_T_1275 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1340 & ~(_T_1275 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1357 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1357 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1357 & ~(_T_1331 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1357 & ~(_T_1331 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1375 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1375 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1375 & ~(_T_1275 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1375 & ~(_T_1275 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1405 & ~(_T_1406 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1405 & ~(_T_1406 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1405 & ~(_T_1410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1405 & ~(_T_1410 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1405 & ~(_T_1414 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1405 & ~(_T_1414 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1405 & ~(_T_1418 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1405 & ~(_T_1418 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1405 & ~(_T_1422 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1405 & ~(_T_1422 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1429 & ~(_T_1430 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1429 & ~(_T_1430 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1429 & ~(_T_1438 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1429 & ~(_T_1438 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1429 & ~(_T_1442 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1429 & ~(_T_1442 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1429 & ~(_T_1450 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1429 & ~(_T_1450 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1459 & ~(_T_1463 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1459 & ~(_T_1463 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1470 & ~(_T_1482 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1470 & ~(_T_1482 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1470 & same_cycle_resp & ~(_T_1488 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1470 & same_cycle_resp & ~(_T_1488 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1470 & same_cycle_resp & ~(_T_1492 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1470 & same_cycle_resp & ~(_T_1492 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1470 & ~same_cycle_resp & ~(_T_1500 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1470 & ~same_cycle_resp & ~(_T_1500 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1470 & ~same_cycle_resp & ~(_T_1504 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1470 & ~same_cycle_resp & ~(_T_1504 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1514 & ~(_T_1516 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1514 & ~(_T_1516 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1523 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1523 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1532 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1532 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1558 & ~(_T_1566[0] | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1558 & ~(_T_1566[0] | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1558 & ~(_T_1576 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1558 & ~(_T_1576 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_1601 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:79:80)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_1601 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[6:0];
  _RAND_10 = {1{`RANDOM}};
  denied = _RAND_10[0:0];
  _RAND_11 = {4{`RANDOM}};
  inflight = _RAND_11[127:0];
  _RAND_12 = {16{`RANDOM}};
  inflight_opcodes = _RAND_12[511:0];
  _RAND_13 = {16{`RANDOM}};
  inflight_sizes = _RAND_13[511:0];
  _RAND_14 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  watchdog = _RAND_16[31:0];
  _RAND_17 = {4{`RANDOM}};
  inflight_1 = _RAND_17[127:0];
  _RAND_18 = {16{`RANDOM}};
  inflight_sizes_1 = _RAND_18[511:0];
  _RAND_19 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  watchdog_1 = _RAND_20[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_17(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [4:0]  io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_echo_tl_state_size,
  input  [6:0]  io_enq_bits_echo_tl_state_source,
  input         io_enq_bits_wen,
  input         io_deq_ready,
  output        io_deq_valid,
  output [4:0]  io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [3:0]  io_deq_bits_echo_tl_state_size,
  output [6:0]  io_deq_bits_echo_tl_state_source,
  output        io_deq_bits_wen
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] ram_id [0:0]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_len [0:0]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_burst [0:0]; // @[Decoupled.scala 218:16]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] ram_echo_tl_state_size [0:0]; // @[Decoupled.scala 218:16]
  wire [3:0] ram_echo_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_echo_tl_state_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [3:0] ram_echo_tl_state_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_echo_tl_state_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_echo_tl_state_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_echo_tl_state_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_echo_tl_state_source [0:0]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_wen [0:0]; // @[Decoupled.scala 218:16]
  wire  ram_wen_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_wen_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_wen_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_wen_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_wen_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_wen_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 249:27 Decoupled.scala 249:36]
  wire  do_enq = empty ? _GEN_18 : _do_enq_T; // @[Decoupled.scala 246:18]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 246:18 Decoupled.scala 248:14]
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_burst_MPORT_data = 2'h1;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_echo_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_size_io_deq_bits_MPORT_data =
    ram_echo_tl_state_size[ram_echo_tl_state_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_echo_tl_state_size_MPORT_data = io_enq_bits_echo_tl_state_size;
  assign ram_echo_tl_state_size_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_size_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_size_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_wen_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wen_io_deq_bits_MPORT_data = ram_wen[ram_wen_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_wen_MPORT_data = io_enq_bits_wen;
  assign ram_wen_MPORT_addr = 1'h0;
  assign ram_wen_MPORT_mask = 1'h1;
  assign ram_wen_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 245:25 Decoupled.scala 245:40 Decoupled.scala 240:16]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_burst = empty ? 2'h1 : ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_echo_tl_state_size = empty ? io_enq_bits_echo_tl_state_size :
    ram_echo_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_echo_tl_state_source = empty ? io_enq_bits_echo_tl_state_source :
    ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  assign io_deq_bits_wen = empty ? io_enq_bits_wen : ram_wen_io_deq_bits_MPORT_data; // @[Decoupled.scala 246:18 Decoupled.scala 247:19 Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_echo_tl_state_size_MPORT_en & ram_echo_tl_state_size_MPORT_mask) begin
      ram_echo_tl_state_size[ram_echo_tl_state_size_MPORT_addr] <= ram_echo_tl_state_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_wen_MPORT_en & ram_wen_MPORT_mask) begin
      ram_wen[ram_wen_MPORT_addr] <= ram_wen_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      if (empty) begin // @[Decoupled.scala 246:18]
        if (io_deq_ready) begin // @[Decoupled.scala 249:27]
          maybe_full <= 1'h0; // @[Decoupled.scala 249:36]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_echo_tl_state_size[initvar] = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_echo_tl_state_source[initvar] = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wen[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLToAXI4(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_a_bits_corrupt,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_awready,
  output        auto_out_awvalid,
  output [4:0]  auto_out_awid,
  output [31:0] auto_out_awaddr,
  output [7:0]  auto_out_awlen,
  output [2:0]  auto_out_awsize,
  output [1:0]  auto_out_awburst,
  output [3:0]  auto_out_awecho_tl_state_size,
  output [6:0]  auto_out_awecho_tl_state_source,
  input         auto_out_wready,
  output        auto_out_wvalid,
  output [63:0] auto_out_wdata,
  output [7:0]  auto_out_wstrb,
  output        auto_out_wlast,
  output        auto_out_bready,
  input         auto_out_bvalid,
  input  [4:0]  auto_out_bid,
  input  [1:0]  auto_out_bresp,
  input  [3:0]  auto_out_becho_tl_state_size,
  input  [6:0]  auto_out_becho_tl_state_source,
  input         auto_out_arready,
  output        auto_out_arvalid,
  output [4:0]  auto_out_arid,
  output [31:0] auto_out_araddr,
  output [7:0]  auto_out_arlen,
  output [2:0]  auto_out_arsize,
  output [1:0]  auto_out_arburst,
  output [3:0]  auto_out_arecho_tl_state_size,
  output [6:0]  auto_out_arecho_tl_state_source,
  output        auto_out_rready,
  input         auto_out_rvalid,
  input  [4:0]  auto_out_rid,
  input  [63:0] auto_out_rdata,
  input  [1:0]  auto_out_rresp,
  input  [3:0]  auto_out_recho_tl_state_size,
  input  [6:0]  auto_out_recho_tl_state_source,
  input         auto_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  deq_clock; // @[Decoupled.scala 296:21]
  wire  deq_reset; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] deq_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [7:0] deq_io_enq_bits_strb; // @[Decoupled.scala 296:21]
  wire  deq_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] deq_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [7:0] deq_io_deq_bits_strb; // @[Decoupled.scala 296:21]
  wire  deq_io_deq_bits_last; // @[Decoupled.scala 296:21]
  wire  queue_arw_deq_clock; // @[Decoupled.scala 296:21]
  wire  queue_arw_deq_reset; // @[Decoupled.scala 296:21]
  wire  queue_arw_deq_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  queue_arw_deq_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] queue_arw_deq_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [31:0] queue_arw_deq_io_enq_bits_addr; // @[Decoupled.scala 296:21]
  wire [7:0] queue_arw_deq_io_enq_bits_len; // @[Decoupled.scala 296:21]
  wire [2:0] queue_arw_deq_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [3:0] queue_arw_deq_io_enq_bits_echo_tl_state_size; // @[Decoupled.scala 296:21]
  wire [6:0] queue_arw_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 296:21]
  wire  queue_arw_deq_io_enq_bits_wen; // @[Decoupled.scala 296:21]
  wire  queue_arw_deq_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  queue_arw_deq_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [31:0] queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 296:21]
  wire [7:0] queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 296:21]
  wire [2:0] queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [1:0] queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 296:21]
  wire [3:0] queue_arw_deq_io_deq_bits_echo_tl_state_size; // @[Decoupled.scala 296:21]
  wire [6:0] queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 296:21]
  wire  queue_arw_deq_io_deq_bits_wen; // @[Decoupled.scala 296:21]
  wire  a_isPut = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [4:0] count_7; // @[ToAXI4.scala 254:28]
  wire  idle_6 = count_7 == 5'h0; // @[ToAXI4.scala 256:26]
  reg  write_6; // @[ToAXI4.scala 255:24]
  wire  mismatch_6 = write_6 != a_isPut; // @[ToAXI4.scala 267:50]
  wire  idStall_6 = ~idle_6 & mismatch_6 | count_7 == 5'h10; // @[ToAXI4.scala 268:34]
  reg [4:0] count_6; // @[ToAXI4.scala 254:28]
  wire  idle_5 = count_6 == 5'h0; // @[ToAXI4.scala 256:26]
  reg  write_5; // @[ToAXI4.scala 255:24]
  wire  mismatch_5 = write_5 != a_isPut; // @[ToAXI4.scala 267:50]
  wire  idStall_5 = ~idle_5 & mismatch_5 | count_6 == 5'h10; // @[ToAXI4.scala 268:34]
  reg [4:0] count_5; // @[ToAXI4.scala 254:28]
  wire  idle_4 = count_5 == 5'h0; // @[ToAXI4.scala 256:26]
  reg  write_4; // @[ToAXI4.scala 255:24]
  wire  mismatch_4 = write_4 != a_isPut; // @[ToAXI4.scala 267:50]
  wire  idStall_4 = ~idle_4 & mismatch_4 | count_5 == 5'h10; // @[ToAXI4.scala 268:34]
  reg [4:0] count_4; // @[ToAXI4.scala 254:28]
  wire  idle_3 = count_4 == 5'h0; // @[ToAXI4.scala 256:26]
  reg  write_3; // @[ToAXI4.scala 255:24]
  wire  mismatch_3 = write_3 != a_isPut; // @[ToAXI4.scala 267:50]
  wire  idStall_3 = ~idle_3 & mismatch_3 | count_4 == 5'h10; // @[ToAXI4.scala 268:34]
  reg [4:0] count_3; // @[ToAXI4.scala 254:28]
  wire  idle_2 = count_3 == 5'h0; // @[ToAXI4.scala 256:26]
  reg  write_2; // @[ToAXI4.scala 255:24]
  wire  mismatch_2 = write_2 != a_isPut; // @[ToAXI4.scala 267:50]
  wire  idStall_2 = ~idle_2 & mismatch_2 | count_3 == 5'h10; // @[ToAXI4.scala 268:34]
  reg [4:0] count_2; // @[ToAXI4.scala 254:28]
  wire  idle_1 = count_2 == 5'h0; // @[ToAXI4.scala 256:26]
  reg  write_1; // @[ToAXI4.scala 255:24]
  wire  mismatch_1 = write_1 != a_isPut; // @[ToAXI4.scala 267:50]
  wire  idStall_1 = ~idle_1 & mismatch_1 | count_2 == 5'h10; // @[ToAXI4.scala 268:34]
  reg [4:0] count_1; // @[ToAXI4.scala 254:28]
  wire  idle = count_1 == 5'h0; // @[ToAXI4.scala 256:26]
  reg  write; // @[ToAXI4.scala 255:24]
  wire  mismatch = write != a_isPut; // @[ToAXI4.scala 267:50]
  wire  idStall_0 = ~idle & mismatch | count_1 == 5'h10; // @[ToAXI4.scala 268:34]
  reg  count_23; // @[ToAXI4.scala 254:28]
  wire  idle_22 = ~count_23; // @[ToAXI4.scala 256:26]
  reg  count_22; // @[ToAXI4.scala 254:28]
  wire  idle_21 = ~count_22; // @[ToAXI4.scala 256:26]
  reg  count_21; // @[ToAXI4.scala 254:28]
  wire  idle_20 = ~count_21; // @[ToAXI4.scala 256:26]
  reg  count_20; // @[ToAXI4.scala 254:28]
  wire  idle_19 = ~count_20; // @[ToAXI4.scala 256:26]
  reg  count_19; // @[ToAXI4.scala 254:28]
  wire  idle_18 = ~count_19; // @[ToAXI4.scala 256:26]
  reg  count_18; // @[ToAXI4.scala 254:28]
  wire  idle_17 = ~count_18; // @[ToAXI4.scala 256:26]
  reg  count_17; // @[ToAXI4.scala 254:28]
  wire  idle_16 = ~count_17; // @[ToAXI4.scala 256:26]
  reg  count_16; // @[ToAXI4.scala 254:28]
  wire  idle_15 = ~count_16; // @[ToAXI4.scala 256:26]
  reg  count_15; // @[ToAXI4.scala 254:28]
  wire  idle_14 = ~count_15; // @[ToAXI4.scala 256:26]
  reg  count_14; // @[ToAXI4.scala 254:28]
  wire  idle_13 = ~count_14; // @[ToAXI4.scala 256:26]
  reg  count_13; // @[ToAXI4.scala 254:28]
  wire  idle_12 = ~count_13; // @[ToAXI4.scala 256:26]
  reg  count_12; // @[ToAXI4.scala 254:28]
  wire  idle_11 = ~count_12; // @[ToAXI4.scala 256:26]
  reg  count_11; // @[ToAXI4.scala 254:28]
  wire  idle_10 = ~count_11; // @[ToAXI4.scala 256:26]
  reg  count_10; // @[ToAXI4.scala 254:28]
  wire  idle_9 = ~count_10; // @[ToAXI4.scala 256:26]
  reg  count_9; // @[ToAXI4.scala 254:28]
  wire  idle_8 = ~count_9; // @[ToAXI4.scala 256:26]
  reg  count_8; // @[ToAXI4.scala 254:28]
  wire  idle_7 = ~count_8; // @[ToAXI4.scala 256:26]
  wire  _GEN_131 = 7'h1 == auto_in_a_bits_source ? count_9 : count_8; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_132 = 7'h2 == auto_in_a_bits_source ? count_10 : _GEN_131; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_133 = 7'h3 == auto_in_a_bits_source ? count_11 : _GEN_132; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_134 = 7'h4 == auto_in_a_bits_source ? count_12 : _GEN_133; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_135 = 7'h5 == auto_in_a_bits_source ? count_13 : _GEN_134; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_136 = 7'h6 == auto_in_a_bits_source ? count_14 : _GEN_135; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_137 = 7'h7 == auto_in_a_bits_source ? count_15 : _GEN_136; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_138 = 7'h8 == auto_in_a_bits_source ? count_16 : _GEN_137; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_139 = 7'h9 == auto_in_a_bits_source ? count_17 : _GEN_138; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_140 = 7'ha == auto_in_a_bits_source ? count_18 : _GEN_139; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_141 = 7'hb == auto_in_a_bits_source ? count_19 : _GEN_140; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_142 = 7'hc == auto_in_a_bits_source ? count_20 : _GEN_141; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_143 = 7'hd == auto_in_a_bits_source ? count_21 : _GEN_142; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_144 = 7'he == auto_in_a_bits_source ? count_22 : _GEN_143; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_145 = 7'hf == auto_in_a_bits_source ? count_23 : _GEN_144; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_146 = 7'h10 == auto_in_a_bits_source ? idStall_0 : _GEN_145; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_147 = 7'h11 == auto_in_a_bits_source ? idStall_0 : _GEN_146; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_148 = 7'h12 == auto_in_a_bits_source ? idStall_0 : _GEN_147; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_149 = 7'h13 == auto_in_a_bits_source ? idStall_0 : _GEN_148; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_150 = 7'h14 == auto_in_a_bits_source ? idStall_0 : _GEN_149; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_151 = 7'h15 == auto_in_a_bits_source ? idStall_0 : _GEN_150; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_152 = 7'h16 == auto_in_a_bits_source ? idStall_0 : _GEN_151; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_153 = 7'h17 == auto_in_a_bits_source ? idStall_0 : _GEN_152; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_154 = 7'h18 == auto_in_a_bits_source ? idStall_0 : _GEN_153; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_155 = 7'h19 == auto_in_a_bits_source ? idStall_0 : _GEN_154; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_156 = 7'h1a == auto_in_a_bits_source ? idStall_0 : _GEN_155; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_157 = 7'h1b == auto_in_a_bits_source ? idStall_0 : _GEN_156; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_158 = 7'h1c == auto_in_a_bits_source ? idStall_0 : _GEN_157; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_159 = 7'h1d == auto_in_a_bits_source ? idStall_0 : _GEN_158; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_160 = 7'h1e == auto_in_a_bits_source ? idStall_0 : _GEN_159; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_161 = 7'h1f == auto_in_a_bits_source ? idStall_0 : _GEN_160; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_162 = 7'h20 == auto_in_a_bits_source ? idStall_1 : _GEN_161; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_163 = 7'h21 == auto_in_a_bits_source ? idStall_1 : _GEN_162; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_164 = 7'h22 == auto_in_a_bits_source ? idStall_1 : _GEN_163; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_165 = 7'h23 == auto_in_a_bits_source ? idStall_1 : _GEN_164; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_166 = 7'h24 == auto_in_a_bits_source ? idStall_1 : _GEN_165; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_167 = 7'h25 == auto_in_a_bits_source ? idStall_1 : _GEN_166; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_168 = 7'h26 == auto_in_a_bits_source ? idStall_1 : _GEN_167; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_169 = 7'h27 == auto_in_a_bits_source ? idStall_1 : _GEN_168; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_170 = 7'h28 == auto_in_a_bits_source ? idStall_1 : _GEN_169; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_171 = 7'h29 == auto_in_a_bits_source ? idStall_1 : _GEN_170; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_172 = 7'h2a == auto_in_a_bits_source ? idStall_1 : _GEN_171; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_173 = 7'h2b == auto_in_a_bits_source ? idStall_1 : _GEN_172; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_174 = 7'h2c == auto_in_a_bits_source ? idStall_1 : _GEN_173; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_175 = 7'h2d == auto_in_a_bits_source ? idStall_1 : _GEN_174; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_176 = 7'h2e == auto_in_a_bits_source ? idStall_1 : _GEN_175; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_177 = 7'h2f == auto_in_a_bits_source ? idStall_1 : _GEN_176; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_178 = 7'h30 == auto_in_a_bits_source ? idStall_2 : _GEN_177; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_179 = 7'h31 == auto_in_a_bits_source ? idStall_2 : _GEN_178; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_180 = 7'h32 == auto_in_a_bits_source ? idStall_2 : _GEN_179; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_181 = 7'h33 == auto_in_a_bits_source ? idStall_2 : _GEN_180; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_182 = 7'h34 == auto_in_a_bits_source ? idStall_2 : _GEN_181; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_183 = 7'h35 == auto_in_a_bits_source ? idStall_2 : _GEN_182; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_184 = 7'h36 == auto_in_a_bits_source ? idStall_2 : _GEN_183; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_185 = 7'h37 == auto_in_a_bits_source ? idStall_2 : _GEN_184; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_186 = 7'h38 == auto_in_a_bits_source ? idStall_2 : _GEN_185; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_187 = 7'h39 == auto_in_a_bits_source ? idStall_2 : _GEN_186; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_188 = 7'h3a == auto_in_a_bits_source ? idStall_2 : _GEN_187; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_189 = 7'h3b == auto_in_a_bits_source ? idStall_2 : _GEN_188; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_190 = 7'h3c == auto_in_a_bits_source ? idStall_2 : _GEN_189; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_191 = 7'h3d == auto_in_a_bits_source ? idStall_2 : _GEN_190; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_192 = 7'h3e == auto_in_a_bits_source ? idStall_2 : _GEN_191; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_193 = 7'h3f == auto_in_a_bits_source ? idStall_2 : _GEN_192; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_194 = 7'h40 == auto_in_a_bits_source ? idStall_3 : _GEN_193; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_195 = 7'h41 == auto_in_a_bits_source ? idStall_3 : _GEN_194; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_196 = 7'h42 == auto_in_a_bits_source ? idStall_3 : _GEN_195; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_197 = 7'h43 == auto_in_a_bits_source ? idStall_3 : _GEN_196; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_198 = 7'h44 == auto_in_a_bits_source ? idStall_3 : _GEN_197; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_199 = 7'h45 == auto_in_a_bits_source ? idStall_3 : _GEN_198; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_200 = 7'h46 == auto_in_a_bits_source ? idStall_3 : _GEN_199; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_201 = 7'h47 == auto_in_a_bits_source ? idStall_3 : _GEN_200; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_202 = 7'h48 == auto_in_a_bits_source ? idStall_3 : _GEN_201; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_203 = 7'h49 == auto_in_a_bits_source ? idStall_3 : _GEN_202; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_204 = 7'h4a == auto_in_a_bits_source ? idStall_3 : _GEN_203; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_205 = 7'h4b == auto_in_a_bits_source ? idStall_3 : _GEN_204; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_206 = 7'h4c == auto_in_a_bits_source ? idStall_3 : _GEN_205; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_207 = 7'h4d == auto_in_a_bits_source ? idStall_3 : _GEN_206; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_208 = 7'h4e == auto_in_a_bits_source ? idStall_3 : _GEN_207; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_209 = 7'h4f == auto_in_a_bits_source ? idStall_3 : _GEN_208; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_210 = 7'h50 == auto_in_a_bits_source ? idStall_4 : _GEN_209; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_211 = 7'h51 == auto_in_a_bits_source ? idStall_4 : _GEN_210; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_212 = 7'h52 == auto_in_a_bits_source ? idStall_4 : _GEN_211; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_213 = 7'h53 == auto_in_a_bits_source ? idStall_4 : _GEN_212; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_214 = 7'h54 == auto_in_a_bits_source ? idStall_4 : _GEN_213; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_215 = 7'h55 == auto_in_a_bits_source ? idStall_4 : _GEN_214; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_216 = 7'h56 == auto_in_a_bits_source ? idStall_4 : _GEN_215; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_217 = 7'h57 == auto_in_a_bits_source ? idStall_4 : _GEN_216; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_218 = 7'h58 == auto_in_a_bits_source ? idStall_4 : _GEN_217; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_219 = 7'h59 == auto_in_a_bits_source ? idStall_4 : _GEN_218; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_220 = 7'h5a == auto_in_a_bits_source ? idStall_4 : _GEN_219; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_221 = 7'h5b == auto_in_a_bits_source ? idStall_4 : _GEN_220; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_222 = 7'h5c == auto_in_a_bits_source ? idStall_4 : _GEN_221; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_223 = 7'h5d == auto_in_a_bits_source ? idStall_4 : _GEN_222; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_224 = 7'h5e == auto_in_a_bits_source ? idStall_4 : _GEN_223; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_225 = 7'h5f == auto_in_a_bits_source ? idStall_4 : _GEN_224; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_226 = 7'h60 == auto_in_a_bits_source ? idStall_5 : _GEN_225; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_227 = 7'h61 == auto_in_a_bits_source ? idStall_5 : _GEN_226; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_228 = 7'h62 == auto_in_a_bits_source ? idStall_5 : _GEN_227; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_229 = 7'h63 == auto_in_a_bits_source ? idStall_5 : _GEN_228; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_230 = 7'h64 == auto_in_a_bits_source ? idStall_5 : _GEN_229; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_231 = 7'h65 == auto_in_a_bits_source ? idStall_5 : _GEN_230; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_232 = 7'h66 == auto_in_a_bits_source ? idStall_5 : _GEN_231; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_233 = 7'h67 == auto_in_a_bits_source ? idStall_5 : _GEN_232; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_234 = 7'h68 == auto_in_a_bits_source ? idStall_5 : _GEN_233; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_235 = 7'h69 == auto_in_a_bits_source ? idStall_5 : _GEN_234; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_236 = 7'h6a == auto_in_a_bits_source ? idStall_5 : _GEN_235; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_237 = 7'h6b == auto_in_a_bits_source ? idStall_5 : _GEN_236; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_238 = 7'h6c == auto_in_a_bits_source ? idStall_5 : _GEN_237; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_239 = 7'h6d == auto_in_a_bits_source ? idStall_5 : _GEN_238; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_240 = 7'h6e == auto_in_a_bits_source ? idStall_5 : _GEN_239; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_241 = 7'h6f == auto_in_a_bits_source ? idStall_5 : _GEN_240; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_242 = 7'h70 == auto_in_a_bits_source ? idStall_6 : _GEN_241; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_243 = 7'h71 == auto_in_a_bits_source ? idStall_6 : _GEN_242; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_244 = 7'h72 == auto_in_a_bits_source ? idStall_6 : _GEN_243; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_245 = 7'h73 == auto_in_a_bits_source ? idStall_6 : _GEN_244; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_246 = 7'h74 == auto_in_a_bits_source ? idStall_6 : _GEN_245; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_247 = 7'h75 == auto_in_a_bits_source ? idStall_6 : _GEN_246; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_248 = 7'h76 == auto_in_a_bits_source ? idStall_6 : _GEN_247; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_249 = 7'h77 == auto_in_a_bits_source ? idStall_6 : _GEN_248; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_250 = 7'h78 == auto_in_a_bits_source ? idStall_6 : _GEN_249; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_251 = 7'h79 == auto_in_a_bits_source ? idStall_6 : _GEN_250; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_252 = 7'h7a == auto_in_a_bits_source ? idStall_6 : _GEN_251; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_253 = 7'h7b == auto_in_a_bits_source ? idStall_6 : _GEN_252; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_254 = 7'h7c == auto_in_a_bits_source ? idStall_6 : _GEN_253; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_255 = 7'h7d == auto_in_a_bits_source ? idStall_6 : _GEN_254; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_256 = 7'h7e == auto_in_a_bits_source ? idStall_6 : _GEN_255; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  wire  _GEN_257 = 7'h7f == auto_in_a_bits_source ? idStall_6 : _GEN_256; // @[ToAXI4.scala 195:49 ToAXI4.scala 195:49]
  reg [2:0] counter; // @[Edges.scala 228:27]
  wire  a_first = counter == 3'h0; // @[Edges.scala 230:25]
  wire  stall = _GEN_257 & a_first; // @[ToAXI4.scala 195:49]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[ToAXI4.scala 196:21]
  reg  doneAW; // @[ToAXI4.scala 161:30]
  wire  out_arw_ready = queue_arw_deq_io_enq_ready; // @[ToAXI4.scala 147:25 Decoupled.scala 299:17]
  wire  _bundleIn_0_a_ready_T_1 = doneAW | out_arw_ready; // @[ToAXI4.scala 196:52]
  wire  out_wready = deq_io_enq_ready; // @[ToAXI4.scala 148:23 Decoupled.scala 299:17]
  wire  _bundleIn_0_a_ready_T_3 = a_isPut ? (doneAW | out_arw_ready) & out_wready : out_arw_ready; // @[ToAXI4.scala 196:34]
  wire  bundleIn_0_a_ready = ~stall & _bundleIn_0_a_ready_T_3; // @[ToAXI4.scala 196:28]
  wire  _T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _beats1_decode_T_1 = 13'h3f << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] beats1_decode = _beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire [2:0] beats1 = a_isPut ? beats1_decode : 3'h0; // @[Edges.scala 220:14]
  wire [2:0] counter1 = counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_last = counter == 3'h1 | beats1 == 3'h0; // @[Edges.scala 231:37]
  wire  queue_arw_bits_wen = queue_arw_deq_io_deq_bits_wen; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  queue_arw_valid = queue_arw_deq_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire [4:0] _GEN_3 = 7'h1 == auto_in_a_bits_source ? 5'h8 : 5'h7; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_4 = 7'h2 == auto_in_a_bits_source ? 5'h9 : _GEN_3; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_5 = 7'h3 == auto_in_a_bits_source ? 5'ha : _GEN_4; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_6 = 7'h4 == auto_in_a_bits_source ? 5'hb : _GEN_5; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_7 = 7'h5 == auto_in_a_bits_source ? 5'hc : _GEN_6; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_8 = 7'h6 == auto_in_a_bits_source ? 5'hd : _GEN_7; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_9 = 7'h7 == auto_in_a_bits_source ? 5'he : _GEN_8; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_10 = 7'h8 == auto_in_a_bits_source ? 5'hf : _GEN_9; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_11 = 7'h9 == auto_in_a_bits_source ? 5'h10 : _GEN_10; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_12 = 7'ha == auto_in_a_bits_source ? 5'h11 : _GEN_11; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_13 = 7'hb == auto_in_a_bits_source ? 5'h12 : _GEN_12; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_14 = 7'hc == auto_in_a_bits_source ? 5'h13 : _GEN_13; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_15 = 7'hd == auto_in_a_bits_source ? 5'h14 : _GEN_14; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_16 = 7'he == auto_in_a_bits_source ? 5'h15 : _GEN_15; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_17 = 7'hf == auto_in_a_bits_source ? 5'h16 : _GEN_16; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_18 = 7'h10 == auto_in_a_bits_source ? 5'h0 : _GEN_17; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_19 = 7'h11 == auto_in_a_bits_source ? 5'h0 : _GEN_18; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_20 = 7'h12 == auto_in_a_bits_source ? 5'h0 : _GEN_19; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_21 = 7'h13 == auto_in_a_bits_source ? 5'h0 : _GEN_20; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_22 = 7'h14 == auto_in_a_bits_source ? 5'h0 : _GEN_21; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_23 = 7'h15 == auto_in_a_bits_source ? 5'h0 : _GEN_22; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_24 = 7'h16 == auto_in_a_bits_source ? 5'h0 : _GEN_23; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_25 = 7'h17 == auto_in_a_bits_source ? 5'h0 : _GEN_24; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_26 = 7'h18 == auto_in_a_bits_source ? 5'h0 : _GEN_25; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_27 = 7'h19 == auto_in_a_bits_source ? 5'h0 : _GEN_26; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_28 = 7'h1a == auto_in_a_bits_source ? 5'h0 : _GEN_27; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_29 = 7'h1b == auto_in_a_bits_source ? 5'h0 : _GEN_28; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_30 = 7'h1c == auto_in_a_bits_source ? 5'h0 : _GEN_29; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_31 = 7'h1d == auto_in_a_bits_source ? 5'h0 : _GEN_30; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_32 = 7'h1e == auto_in_a_bits_source ? 5'h0 : _GEN_31; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_33 = 7'h1f == auto_in_a_bits_source ? 5'h0 : _GEN_32; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_34 = 7'h20 == auto_in_a_bits_source ? 5'h1 : _GEN_33; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_35 = 7'h21 == auto_in_a_bits_source ? 5'h1 : _GEN_34; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_36 = 7'h22 == auto_in_a_bits_source ? 5'h1 : _GEN_35; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_37 = 7'h23 == auto_in_a_bits_source ? 5'h1 : _GEN_36; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_38 = 7'h24 == auto_in_a_bits_source ? 5'h1 : _GEN_37; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_39 = 7'h25 == auto_in_a_bits_source ? 5'h1 : _GEN_38; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_40 = 7'h26 == auto_in_a_bits_source ? 5'h1 : _GEN_39; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_41 = 7'h27 == auto_in_a_bits_source ? 5'h1 : _GEN_40; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_42 = 7'h28 == auto_in_a_bits_source ? 5'h1 : _GEN_41; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_43 = 7'h29 == auto_in_a_bits_source ? 5'h1 : _GEN_42; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_44 = 7'h2a == auto_in_a_bits_source ? 5'h1 : _GEN_43; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_45 = 7'h2b == auto_in_a_bits_source ? 5'h1 : _GEN_44; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_46 = 7'h2c == auto_in_a_bits_source ? 5'h1 : _GEN_45; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_47 = 7'h2d == auto_in_a_bits_source ? 5'h1 : _GEN_46; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_48 = 7'h2e == auto_in_a_bits_source ? 5'h1 : _GEN_47; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_49 = 7'h2f == auto_in_a_bits_source ? 5'h1 : _GEN_48; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_50 = 7'h30 == auto_in_a_bits_source ? 5'h2 : _GEN_49; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_51 = 7'h31 == auto_in_a_bits_source ? 5'h2 : _GEN_50; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_52 = 7'h32 == auto_in_a_bits_source ? 5'h2 : _GEN_51; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_53 = 7'h33 == auto_in_a_bits_source ? 5'h2 : _GEN_52; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_54 = 7'h34 == auto_in_a_bits_source ? 5'h2 : _GEN_53; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_55 = 7'h35 == auto_in_a_bits_source ? 5'h2 : _GEN_54; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_56 = 7'h36 == auto_in_a_bits_source ? 5'h2 : _GEN_55; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_57 = 7'h37 == auto_in_a_bits_source ? 5'h2 : _GEN_56; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_58 = 7'h38 == auto_in_a_bits_source ? 5'h2 : _GEN_57; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_59 = 7'h39 == auto_in_a_bits_source ? 5'h2 : _GEN_58; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_60 = 7'h3a == auto_in_a_bits_source ? 5'h2 : _GEN_59; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_61 = 7'h3b == auto_in_a_bits_source ? 5'h2 : _GEN_60; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_62 = 7'h3c == auto_in_a_bits_source ? 5'h2 : _GEN_61; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_63 = 7'h3d == auto_in_a_bits_source ? 5'h2 : _GEN_62; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_64 = 7'h3e == auto_in_a_bits_source ? 5'h2 : _GEN_63; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_65 = 7'h3f == auto_in_a_bits_source ? 5'h2 : _GEN_64; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_66 = 7'h40 == auto_in_a_bits_source ? 5'h3 : _GEN_65; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_67 = 7'h41 == auto_in_a_bits_source ? 5'h3 : _GEN_66; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_68 = 7'h42 == auto_in_a_bits_source ? 5'h3 : _GEN_67; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_69 = 7'h43 == auto_in_a_bits_source ? 5'h3 : _GEN_68; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_70 = 7'h44 == auto_in_a_bits_source ? 5'h3 : _GEN_69; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_71 = 7'h45 == auto_in_a_bits_source ? 5'h3 : _GEN_70; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_72 = 7'h46 == auto_in_a_bits_source ? 5'h3 : _GEN_71; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_73 = 7'h47 == auto_in_a_bits_source ? 5'h3 : _GEN_72; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_74 = 7'h48 == auto_in_a_bits_source ? 5'h3 : _GEN_73; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_75 = 7'h49 == auto_in_a_bits_source ? 5'h3 : _GEN_74; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_76 = 7'h4a == auto_in_a_bits_source ? 5'h3 : _GEN_75; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_77 = 7'h4b == auto_in_a_bits_source ? 5'h3 : _GEN_76; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_78 = 7'h4c == auto_in_a_bits_source ? 5'h3 : _GEN_77; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_79 = 7'h4d == auto_in_a_bits_source ? 5'h3 : _GEN_78; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_80 = 7'h4e == auto_in_a_bits_source ? 5'h3 : _GEN_79; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_81 = 7'h4f == auto_in_a_bits_source ? 5'h3 : _GEN_80; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_82 = 7'h50 == auto_in_a_bits_source ? 5'h4 : _GEN_81; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_83 = 7'h51 == auto_in_a_bits_source ? 5'h4 : _GEN_82; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_84 = 7'h52 == auto_in_a_bits_source ? 5'h4 : _GEN_83; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_85 = 7'h53 == auto_in_a_bits_source ? 5'h4 : _GEN_84; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_86 = 7'h54 == auto_in_a_bits_source ? 5'h4 : _GEN_85; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_87 = 7'h55 == auto_in_a_bits_source ? 5'h4 : _GEN_86; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_88 = 7'h56 == auto_in_a_bits_source ? 5'h4 : _GEN_87; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_89 = 7'h57 == auto_in_a_bits_source ? 5'h4 : _GEN_88; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_90 = 7'h58 == auto_in_a_bits_source ? 5'h4 : _GEN_89; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_91 = 7'h59 == auto_in_a_bits_source ? 5'h4 : _GEN_90; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_92 = 7'h5a == auto_in_a_bits_source ? 5'h4 : _GEN_91; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_93 = 7'h5b == auto_in_a_bits_source ? 5'h4 : _GEN_92; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_94 = 7'h5c == auto_in_a_bits_source ? 5'h4 : _GEN_93; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_95 = 7'h5d == auto_in_a_bits_source ? 5'h4 : _GEN_94; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_96 = 7'h5e == auto_in_a_bits_source ? 5'h4 : _GEN_95; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_97 = 7'h5f == auto_in_a_bits_source ? 5'h4 : _GEN_96; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_98 = 7'h60 == auto_in_a_bits_source ? 5'h5 : _GEN_97; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_99 = 7'h61 == auto_in_a_bits_source ? 5'h5 : _GEN_98; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_100 = 7'h62 == auto_in_a_bits_source ? 5'h5 : _GEN_99; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_101 = 7'h63 == auto_in_a_bits_source ? 5'h5 : _GEN_100; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_102 = 7'h64 == auto_in_a_bits_source ? 5'h5 : _GEN_101; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_103 = 7'h65 == auto_in_a_bits_source ? 5'h5 : _GEN_102; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_104 = 7'h66 == auto_in_a_bits_source ? 5'h5 : _GEN_103; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_105 = 7'h67 == auto_in_a_bits_source ? 5'h5 : _GEN_104; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_106 = 7'h68 == auto_in_a_bits_source ? 5'h5 : _GEN_105; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_107 = 7'h69 == auto_in_a_bits_source ? 5'h5 : _GEN_106; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_108 = 7'h6a == auto_in_a_bits_source ? 5'h5 : _GEN_107; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_109 = 7'h6b == auto_in_a_bits_source ? 5'h5 : _GEN_108; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_110 = 7'h6c == auto_in_a_bits_source ? 5'h5 : _GEN_109; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_111 = 7'h6d == auto_in_a_bits_source ? 5'h5 : _GEN_110; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_112 = 7'h6e == auto_in_a_bits_source ? 5'h5 : _GEN_111; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_113 = 7'h6f == auto_in_a_bits_source ? 5'h5 : _GEN_112; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_114 = 7'h70 == auto_in_a_bits_source ? 5'h6 : _GEN_113; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_115 = 7'h71 == auto_in_a_bits_source ? 5'h6 : _GEN_114; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_116 = 7'h72 == auto_in_a_bits_source ? 5'h6 : _GEN_115; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_117 = 7'h73 == auto_in_a_bits_source ? 5'h6 : _GEN_116; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_118 = 7'h74 == auto_in_a_bits_source ? 5'h6 : _GEN_117; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_119 = 7'h75 == auto_in_a_bits_source ? 5'h6 : _GEN_118; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_120 = 7'h76 == auto_in_a_bits_source ? 5'h6 : _GEN_119; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_121 = 7'h77 == auto_in_a_bits_source ? 5'h6 : _GEN_120; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_122 = 7'h78 == auto_in_a_bits_source ? 5'h6 : _GEN_121; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_123 = 7'h79 == auto_in_a_bits_source ? 5'h6 : _GEN_122; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_124 = 7'h7a == auto_in_a_bits_source ? 5'h6 : _GEN_123; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_125 = 7'h7b == auto_in_a_bits_source ? 5'h6 : _GEN_124; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_126 = 7'h7c == auto_in_a_bits_source ? 5'h6 : _GEN_125; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_127 = 7'h7d == auto_in_a_bits_source ? 5'h6 : _GEN_126; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] _GEN_128 = 7'h7e == auto_in_a_bits_source ? 5'h6 : _GEN_127; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [4:0] out_arw_bits_id = 7'h7f == auto_in_a_bits_source ? 5'h6 : _GEN_128; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  wire [17:0] _out_arw_bits_len_T_1 = 18'h7ff << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [10:0] _out_arw_bits_len_T_3 = ~_out_arw_bits_len_T_1[10:0]; // @[package.scala 234:46]
  wire  _out_arw_valid_T_1 = _bundleIn_0_a_ready_T & auto_in_a_valid; // @[ToAXI4.scala 197:31]
  wire  _out_arw_valid_T_4 = a_isPut ? ~doneAW & out_wready : 1'h1; // @[ToAXI4.scala 197:51]
  wire  out_arw_valid = _bundleIn_0_a_ready_T & auto_in_a_valid & _out_arw_valid_T_4; // @[ToAXI4.scala 197:45]
  reg  r_holds_d; // @[ToAXI4.scala 206:30]
  reg [2:0] b_delay; // @[ToAXI4.scala 209:24]
  wire  r_wins = auto_out_rvalid & b_delay != 3'h7 | r_holds_d; // @[ToAXI4.scala 215:57]
  wire  bundleOut_0_rready = auto_in_d_ready & r_wins; // @[ToAXI4.scala 217:33]
  wire  _T_2 = bundleOut_0_rready & auto_out_rvalid; // @[Decoupled.scala 40:37]
  wire  bundleOut_0_bready = auto_in_d_ready & ~r_wins; // @[ToAXI4.scala 218:33]
  wire [2:0] _bdelay_T_1 = b_delay + 3'h1; // @[ToAXI4.scala 211:28]
  wire  bundleIn_0_d_valid = r_wins ? auto_out_rvalid : auto_out_bvalid; // @[ToAXI4.scala 219:24]
  reg  r_first; // @[ToAXI4.scala 224:28]
  wire  _GEN_260 = _T_2 ? auto_out_rlast : r_first; // @[ToAXI4.scala 225:27 ToAXI4.scala 225:37 ToAXI4.scala 224:28]
  wire  _rdenied_T = auto_out_rresp == 2'h3; // @[ToAXI4.scala 226:39]
  reg  r_denied_r; // @[Reg.scala 15:16]
  wire  _GEN_261 = r_first ? _rdenied_T : r_denied_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire  r_corrupt = auto_out_rresp != 2'h0; // @[ToAXI4.scala 227:39]
  wire  b_denied = auto_out_bresp != 2'h0; // @[ToAXI4.scala 228:39]
  wire  r_d_corrupt = r_corrupt | _GEN_261; // @[ToAXI4.scala 230:100]
  wire [2:0] r_d_size = auto_out_recho_tl_state_size[2:0]; // @[Edges.scala 771:17 Edges.scala 774:15]
  wire [2:0] b_d_size = auto_out_becho_tl_state_size[2:0]; // @[Edges.scala 755:17 Edges.scala 758:15]
  wire [31:0] _a_sel_T = 32'h1 << out_arw_bits_id; // @[OneHot.scala 65:12]
  wire  a_sel_0 = _a_sel_T[0]; // @[ToAXI4.scala 242:58]
  wire  a_sel_1 = _a_sel_T[1]; // @[ToAXI4.scala 242:58]
  wire  a_sel_2 = _a_sel_T[2]; // @[ToAXI4.scala 242:58]
  wire  a_sel_3 = _a_sel_T[3]; // @[ToAXI4.scala 242:58]
  wire  a_sel_4 = _a_sel_T[4]; // @[ToAXI4.scala 242:58]
  wire  a_sel_5 = _a_sel_T[5]; // @[ToAXI4.scala 242:58]
  wire  a_sel_6 = _a_sel_T[6]; // @[ToAXI4.scala 242:58]
  wire  a_sel_7 = _a_sel_T[7]; // @[ToAXI4.scala 242:58]
  wire  a_sel_8 = _a_sel_T[8]; // @[ToAXI4.scala 242:58]
  wire  a_sel_9 = _a_sel_T[9]; // @[ToAXI4.scala 242:58]
  wire  a_sel_10 = _a_sel_T[10]; // @[ToAXI4.scala 242:58]
  wire  a_sel_11 = _a_sel_T[11]; // @[ToAXI4.scala 242:58]
  wire  a_sel_12 = _a_sel_T[12]; // @[ToAXI4.scala 242:58]
  wire  a_sel_13 = _a_sel_T[13]; // @[ToAXI4.scala 242:58]
  wire  a_sel_14 = _a_sel_T[14]; // @[ToAXI4.scala 242:58]
  wire  a_sel_15 = _a_sel_T[15]; // @[ToAXI4.scala 242:58]
  wire  a_sel_16 = _a_sel_T[16]; // @[ToAXI4.scala 242:58]
  wire  a_sel_17 = _a_sel_T[17]; // @[ToAXI4.scala 242:58]
  wire  a_sel_18 = _a_sel_T[18]; // @[ToAXI4.scala 242:58]
  wire  a_sel_19 = _a_sel_T[19]; // @[ToAXI4.scala 242:58]
  wire  a_sel_20 = _a_sel_T[20]; // @[ToAXI4.scala 242:58]
  wire  a_sel_21 = _a_sel_T[21]; // @[ToAXI4.scala 242:58]
  wire  a_sel_22 = _a_sel_T[22]; // @[ToAXI4.scala 242:58]
  wire [4:0] d_sel_shiftAmount = r_wins ? auto_out_rid : auto_out_bid; // @[ToAXI4.scala 243:31]
  wire [31:0] _d_sel_T_1 = 32'h1 << d_sel_shiftAmount; // @[OneHot.scala 65:12]
  wire  d_sel_0 = _d_sel_T_1[0]; // @[ToAXI4.scala 243:93]
  wire  d_sel_1 = _d_sel_T_1[1]; // @[ToAXI4.scala 243:93]
  wire  d_sel_2 = _d_sel_T_1[2]; // @[ToAXI4.scala 243:93]
  wire  d_sel_3 = _d_sel_T_1[3]; // @[ToAXI4.scala 243:93]
  wire  d_sel_4 = _d_sel_T_1[4]; // @[ToAXI4.scala 243:93]
  wire  d_sel_5 = _d_sel_T_1[5]; // @[ToAXI4.scala 243:93]
  wire  d_sel_6 = _d_sel_T_1[6]; // @[ToAXI4.scala 243:93]
  wire  d_sel_7 = _d_sel_T_1[7]; // @[ToAXI4.scala 243:93]
  wire  d_sel_8 = _d_sel_T_1[8]; // @[ToAXI4.scala 243:93]
  wire  d_sel_9 = _d_sel_T_1[9]; // @[ToAXI4.scala 243:93]
  wire  d_sel_10 = _d_sel_T_1[10]; // @[ToAXI4.scala 243:93]
  wire  d_sel_11 = _d_sel_T_1[11]; // @[ToAXI4.scala 243:93]
  wire  d_sel_12 = _d_sel_T_1[12]; // @[ToAXI4.scala 243:93]
  wire  d_sel_13 = _d_sel_T_1[13]; // @[ToAXI4.scala 243:93]
  wire  d_sel_14 = _d_sel_T_1[14]; // @[ToAXI4.scala 243:93]
  wire  d_sel_15 = _d_sel_T_1[15]; // @[ToAXI4.scala 243:93]
  wire  d_sel_16 = _d_sel_T_1[16]; // @[ToAXI4.scala 243:93]
  wire  d_sel_17 = _d_sel_T_1[17]; // @[ToAXI4.scala 243:93]
  wire  d_sel_18 = _d_sel_T_1[18]; // @[ToAXI4.scala 243:93]
  wire  d_sel_19 = _d_sel_T_1[19]; // @[ToAXI4.scala 243:93]
  wire  d_sel_20 = _d_sel_T_1[20]; // @[ToAXI4.scala 243:93]
  wire  d_sel_21 = _d_sel_T_1[21]; // @[ToAXI4.scala 243:93]
  wire  d_sel_22 = _d_sel_T_1[22]; // @[ToAXI4.scala 243:93]
  wire  d_last = r_wins ? auto_out_rlast : 1'h1; // @[ToAXI4.scala 244:23]
  wire  _inc_T = out_arw_ready & out_arw_valid; // @[Decoupled.scala 40:37]
  wire  inc = a_sel_0 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  _dec_T_1 = auto_in_d_ready & bundleIn_0_d_valid; // @[Decoupled.scala 40:37]
  wire  dec = d_sel_0 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire [4:0] _GEN_285 = {{4'd0}, inc}; // @[ToAXI4.scala 260:24]
  wire [4:0] _count_T_2 = count_1 + _GEN_285; // @[ToAXI4.scala 260:24]
  wire [4:0] _GEN_286 = {{4'd0}, dec}; // @[ToAXI4.scala 260:37]
  wire [4:0] _count_T_4 = _count_T_2 - _GEN_286; // @[ToAXI4.scala 260:37]
  wire  inc_1 = a_sel_1 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_1 = d_sel_1 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire [4:0] _GEN_287 = {{4'd0}, inc_1}; // @[ToAXI4.scala 260:24]
  wire [4:0] _count_T_6 = count_2 + _GEN_287; // @[ToAXI4.scala 260:24]
  wire [4:0] _GEN_288 = {{4'd0}, dec_1}; // @[ToAXI4.scala 260:37]
  wire [4:0] _count_T_8 = _count_T_6 - _GEN_288; // @[ToAXI4.scala 260:37]
  wire  inc_2 = a_sel_2 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_2 = d_sel_2 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire [4:0] _GEN_289 = {{4'd0}, inc_2}; // @[ToAXI4.scala 260:24]
  wire [4:0] _count_T_10 = count_3 + _GEN_289; // @[ToAXI4.scala 260:24]
  wire [4:0] _GEN_290 = {{4'd0}, dec_2}; // @[ToAXI4.scala 260:37]
  wire [4:0] _count_T_12 = _count_T_10 - _GEN_290; // @[ToAXI4.scala 260:37]
  wire  inc_3 = a_sel_3 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_3 = d_sel_3 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire [4:0] _GEN_291 = {{4'd0}, inc_3}; // @[ToAXI4.scala 260:24]
  wire [4:0] _count_T_14 = count_4 + _GEN_291; // @[ToAXI4.scala 260:24]
  wire [4:0] _GEN_292 = {{4'd0}, dec_3}; // @[ToAXI4.scala 260:37]
  wire [4:0] _count_T_16 = _count_T_14 - _GEN_292; // @[ToAXI4.scala 260:37]
  wire  inc_4 = a_sel_4 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_4 = d_sel_4 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire [4:0] _GEN_293 = {{4'd0}, inc_4}; // @[ToAXI4.scala 260:24]
  wire [4:0] _count_T_18 = count_5 + _GEN_293; // @[ToAXI4.scala 260:24]
  wire [4:0] _GEN_294 = {{4'd0}, dec_4}; // @[ToAXI4.scala 260:37]
  wire [4:0] _count_T_20 = _count_T_18 - _GEN_294; // @[ToAXI4.scala 260:37]
  wire  inc_5 = a_sel_5 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_5 = d_sel_5 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire [4:0] _GEN_295 = {{4'd0}, inc_5}; // @[ToAXI4.scala 260:24]
  wire [4:0] _count_T_22 = count_6 + _GEN_295; // @[ToAXI4.scala 260:24]
  wire [4:0] _GEN_296 = {{4'd0}, dec_5}; // @[ToAXI4.scala 260:37]
  wire [4:0] _count_T_24 = _count_T_22 - _GEN_296; // @[ToAXI4.scala 260:37]
  wire  inc_6 = a_sel_6 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_6 = d_sel_6 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire [4:0] _GEN_297 = {{4'd0}, inc_6}; // @[ToAXI4.scala 260:24]
  wire [4:0] _count_T_26 = count_7 + _GEN_297; // @[ToAXI4.scala 260:24]
  wire [4:0] _GEN_298 = {{4'd0}, dec_6}; // @[ToAXI4.scala 260:37]
  wire [4:0] _count_T_28 = _count_T_26 - _GEN_298; // @[ToAXI4.scala 260:37]
  wire  inc_7 = a_sel_7 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_7 = d_sel_7 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_30 = count_8 + inc_7; // @[ToAXI4.scala 260:24]
  wire  inc_8 = a_sel_8 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_8 = d_sel_8 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_34 = count_9 + inc_8; // @[ToAXI4.scala 260:24]
  wire  inc_9 = a_sel_9 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_9 = d_sel_9 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_38 = count_10 + inc_9; // @[ToAXI4.scala 260:24]
  wire  inc_10 = a_sel_10 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_10 = d_sel_10 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_42 = count_11 + inc_10; // @[ToAXI4.scala 260:24]
  wire  inc_11 = a_sel_11 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_11 = d_sel_11 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_46 = count_12 + inc_11; // @[ToAXI4.scala 260:24]
  wire  inc_12 = a_sel_12 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_12 = d_sel_12 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_50 = count_13 + inc_12; // @[ToAXI4.scala 260:24]
  wire  inc_13 = a_sel_13 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_13 = d_sel_13 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_54 = count_14 + inc_13; // @[ToAXI4.scala 260:24]
  wire  inc_14 = a_sel_14 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_14 = d_sel_14 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_58 = count_15 + inc_14; // @[ToAXI4.scala 260:24]
  wire  inc_15 = a_sel_15 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_15 = d_sel_15 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_62 = count_16 + inc_15; // @[ToAXI4.scala 260:24]
  wire  inc_16 = a_sel_16 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_16 = d_sel_16 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_66 = count_17 + inc_16; // @[ToAXI4.scala 260:24]
  wire  inc_17 = a_sel_17 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_17 = d_sel_17 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_70 = count_18 + inc_17; // @[ToAXI4.scala 260:24]
  wire  inc_18 = a_sel_18 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_18 = d_sel_18 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_74 = count_19 + inc_18; // @[ToAXI4.scala 260:24]
  wire  inc_19 = a_sel_19 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_19 = d_sel_19 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_78 = count_20 + inc_19; // @[ToAXI4.scala 260:24]
  wire  inc_20 = a_sel_20 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_20 = d_sel_20 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_82 = count_21 + inc_20; // @[ToAXI4.scala 260:24]
  wire  inc_21 = a_sel_21 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_21 = d_sel_21 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_86 = count_22 + inc_21; // @[ToAXI4.scala 260:24]
  wire  inc_22 = a_sel_22 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_22 = d_sel_22 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _count_T_90 = count_23 + inc_22; // @[ToAXI4.scala 260:24]
  TLMonitor_10 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_15 deq ( // @[Decoupled.scala 296:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_data(deq_io_enq_bits_data),
    .io_enq_bits_strb(deq_io_enq_bits_strb),
    .io_enq_bits_last(deq_io_enq_bits_last),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_data(deq_io_deq_bits_data),
    .io_deq_bits_strb(deq_io_deq_bits_strb),
    .io_deq_bits_last(deq_io_deq_bits_last)
  );
  Queue_17 queue_arw_deq ( // @[Decoupled.scala 296:21]
    .clock(queue_arw_deq_clock),
    .reset(queue_arw_deq_reset),
    .io_enq_ready(queue_arw_deq_io_enq_ready),
    .io_enq_valid(queue_arw_deq_io_enq_valid),
    .io_enq_bits_id(queue_arw_deq_io_enq_bits_id),
    .io_enq_bits_addr(queue_arw_deq_io_enq_bits_addr),
    .io_enq_bits_len(queue_arw_deq_io_enq_bits_len),
    .io_enq_bits_size(queue_arw_deq_io_enq_bits_size),
    .io_enq_bits_echo_tl_state_size(queue_arw_deq_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(queue_arw_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_wen(queue_arw_deq_io_enq_bits_wen),
    .io_deq_ready(queue_arw_deq_io_deq_ready),
    .io_deq_valid(queue_arw_deq_io_deq_valid),
    .io_deq_bits_id(queue_arw_deq_io_deq_bits_id),
    .io_deq_bits_addr(queue_arw_deq_io_deq_bits_addr),
    .io_deq_bits_len(queue_arw_deq_io_deq_bits_len),
    .io_deq_bits_size(queue_arw_deq_io_deq_bits_size),
    .io_deq_bits_burst(queue_arw_deq_io_deq_bits_burst),
    .io_deq_bits_echo_tl_state_size(queue_arw_deq_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(queue_arw_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_wen(queue_arw_deq_io_deq_bits_wen)
  );
  assign auto_in_a_ready = ~stall & _bundleIn_0_a_ready_T_3; // @[ToAXI4.scala 196:28]
  assign auto_in_d_valid = r_wins ? auto_out_rvalid : auto_out_bvalid; // @[ToAXI4.scala 219:24]
  assign auto_in_d_bits_opcode = r_wins ? 3'h1 : 3'h0; // @[ToAXI4.scala 237:23]
  assign auto_in_d_bits_size = r_wins ? r_d_size : b_d_size; // @[ToAXI4.scala 237:23]
  assign auto_in_d_bits_source = r_wins ? auto_out_recho_tl_state_source : auto_out_becho_tl_state_source; // @[ToAXI4.scala 237:23]
  assign auto_in_d_bits_denied = r_wins ? _GEN_261 : b_denied; // @[ToAXI4.scala 237:23]
  assign auto_in_d_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = r_wins & r_d_corrupt; // @[ToAXI4.scala 237:23]
  assign auto_out_awvalid = queue_arw_valid & queue_arw_bits_wen; // @[ToAXI4.scala 156:39]
  assign auto_out_awid = queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awaddr = queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awlen = queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awsize = queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awburst = queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awecho_tl_state_size = queue_arw_deq_io_deq_bits_echo_tl_state_size; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_awecho_tl_state_source = queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_wvalid = deq_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  assign auto_out_wdata = deq_io_deq_bits_data; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_wstrb = deq_io_deq_bits_strb; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_wlast = deq_io_deq_bits_last; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_bready = auto_in_d_ready & ~r_wins; // @[ToAXI4.scala 218:33]
  assign auto_out_arvalid = queue_arw_valid & ~queue_arw_bits_wen; // @[ToAXI4.scala 155:39]
  assign auto_out_arid = queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_araddr = queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_arlen = queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_arsize = queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_arburst = queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_arecho_tl_state_size = queue_arw_deq_io_deq_bits_echo_tl_state_size; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_arecho_tl_state_source = queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  assign auto_out_rready = auto_in_d_ready & r_wins; // @[ToAXI4.scala 217:33]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = ~stall & _bundleIn_0_a_ready_T_3; // @[ToAXI4.scala 196:28]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = r_wins ? auto_out_rvalid : auto_out_bvalid; // @[ToAXI4.scala 219:24]
  assign monitor_io_in_d_bits_opcode = r_wins ? 3'h1 : 3'h0; // @[ToAXI4.scala 237:23]
  assign monitor_io_in_d_bits_size = r_wins ? r_d_size : b_d_size; // @[ToAXI4.scala 237:23]
  assign monitor_io_in_d_bits_source = r_wins ? auto_out_recho_tl_state_source :
    auto_out_becho_tl_state_source; // @[ToAXI4.scala 237:23]
  assign monitor_io_in_d_bits_denied = r_wins ? _GEN_261 : b_denied; // @[ToAXI4.scala 237:23]
  assign monitor_io_in_d_bits_corrupt = r_wins & r_d_corrupt; // @[ToAXI4.scala 237:23]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = _out_arw_valid_T_1 & a_isPut & _bundleIn_0_a_ready_T_1; // @[ToAXI4.scala 199:54]
  assign deq_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_strb = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_last = counter == 3'h1 | beats1 == 3'h0; // @[Edges.scala 231:37]
  assign deq_io_deq_ready = auto_out_wready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign queue_arw_deq_clock = clock;
  assign queue_arw_deq_reset = reset;
  assign queue_arw_deq_io_enq_valid = _bundleIn_0_a_ready_T & auto_in_a_valid & _out_arw_valid_T_4; // @[ToAXI4.scala 197:45]
  assign queue_arw_deq_io_enq_bits_id = 7'h7f == auto_in_a_bits_source ? 5'h6 : _GEN_128; // @[ToAXI4.scala 166:17 ToAXI4.scala 166:17]
  assign queue_arw_deq_io_enq_bits_addr = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign queue_arw_deq_io_enq_bits_len = _out_arw_bits_len_T_3[10:3]; // @[ToAXI4.scala 168:84]
  assign queue_arw_deq_io_enq_bits_size = auto_in_a_bits_size >= 3'h3 ? 3'h3 : auto_in_a_bits_size; // @[ToAXI4.scala 169:23]
  assign queue_arw_deq_io_enq_bits_echo_tl_state_size = {{1'd0}, auto_in_a_bits_size}; // @[ToAXI4.scala 147:25 ToAXI4.scala 179:22]
  assign queue_arw_deq_io_enq_bits_echo_tl_state_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign queue_arw_deq_io_enq_bits_wen = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  assign queue_arw_deq_io_deq_ready = queue_arw_bits_wen ? auto_out_awready : auto_out_arready; // @[ToAXI4.scala 157:29]
  always @(posedge clock) begin
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_7 <= 5'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_7 <= _count_T_28; // @[ToAXI4.scala 260:15]
    end
    if (inc_6) begin // @[ToAXI4.scala 265:20]
      write_6 <= a_isPut; // @[ToAXI4.scala 265:28]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_6 <= 5'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_6 <= _count_T_24; // @[ToAXI4.scala 260:15]
    end
    if (inc_5) begin // @[ToAXI4.scala 265:20]
      write_5 <= a_isPut; // @[ToAXI4.scala 265:28]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_5 <= 5'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_5 <= _count_T_20; // @[ToAXI4.scala 260:15]
    end
    if (inc_4) begin // @[ToAXI4.scala 265:20]
      write_4 <= a_isPut; // @[ToAXI4.scala 265:28]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_4 <= 5'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_4 <= _count_T_16; // @[ToAXI4.scala 260:15]
    end
    if (inc_3) begin // @[ToAXI4.scala 265:20]
      write_3 <= a_isPut; // @[ToAXI4.scala 265:28]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_3 <= 5'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_3 <= _count_T_12; // @[ToAXI4.scala 260:15]
    end
    if (inc_2) begin // @[ToAXI4.scala 265:20]
      write_2 <= a_isPut; // @[ToAXI4.scala 265:28]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_2 <= 5'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_2 <= _count_T_8; // @[ToAXI4.scala 260:15]
    end
    if (inc_1) begin // @[ToAXI4.scala 265:20]
      write_1 <= a_isPut; // @[ToAXI4.scala 265:28]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_1 <= 5'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_1 <= _count_T_4; // @[ToAXI4.scala 260:15]
    end
    if (inc) begin // @[ToAXI4.scala 265:20]
      write <= a_isPut; // @[ToAXI4.scala 265:28]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_23 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_23 <= _count_T_90 - dec_22; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_22 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_22 <= _count_T_86 - dec_21; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_21 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_21 <= _count_T_82 - dec_20; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_20 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_20 <= _count_T_78 - dec_19; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_19 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_19 <= _count_T_74 - dec_18; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_18 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_18 <= _count_T_70 - dec_17; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_17 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_17 <= _count_T_66 - dec_16; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_16 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_16 <= _count_T_62 - dec_15; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_15 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_15 <= _count_T_58 - dec_14; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_14 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_14 <= _count_T_54 - dec_13; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_13 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_13 <= _count_T_50 - dec_12; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_12 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_12 <= _count_T_46 - dec_11; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_11 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_11 <= _count_T_42 - dec_10; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_10 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_10 <= _count_T_38 - dec_9; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_9 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_9 <= _count_T_34 - dec_8; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_8 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_8 <= _count_T_30 - dec_7; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_isPut) begin // @[Edges.scala 220:14]
          counter <= beats1_decode;
        end else begin
          counter <= 3'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (reset) begin // @[ToAXI4.scala 161:30]
      doneAW <= 1'h0; // @[ToAXI4.scala 161:30]
    end else if (_T) begin // @[ToAXI4.scala 162:26]
      doneAW <= ~a_last; // @[ToAXI4.scala 162:35]
    end
    if (reset) begin // @[ToAXI4.scala 206:30]
      r_holds_d <= 1'h0; // @[ToAXI4.scala 206:30]
    end else if (_T_2) begin // @[ToAXI4.scala 207:27]
      r_holds_d <= ~auto_out_rlast; // @[ToAXI4.scala 207:39]
    end
    if (auto_out_bvalid & ~bundleOut_0_bready) begin // @[ToAXI4.scala 210:42]
      b_delay <= _bdelay_T_1; // @[ToAXI4.scala 211:17]
    end else begin
      b_delay <= 3'h0; // @[ToAXI4.scala 213:17]
    end
    r_first <= reset | _GEN_260; // @[ToAXI4.scala 224:28 ToAXI4.scala 224:28]
    if (r_first) begin // @[Reg.scala 16:19]
      r_denied_r <= _rdenied_T; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec | count_1 != 5'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec | count_1 != 5'h0 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc | count_1 != 5'h10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc | count_1 != 5'h10 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_1 | count_2 != 5'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_1 | count_2 != 5'h0 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_1 | count_2 != 5'h10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_1 | count_2 != 5'h10 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_2 | count_3 != 5'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_2 | count_3 != 5'h0 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_2 | count_3 != 5'h10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_2 | count_3 != 5'h10 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_3 | count_4 != 5'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_3 | count_4 != 5'h0 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_3 | count_4 != 5'h10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_3 | count_4 != 5'h10 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_4 | count_5 != 5'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_4 | count_5 != 5'h0 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_4 | count_5 != 5'h10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_4 | count_5 != 5'h10 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_5 | count_6 != 5'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_5 | count_6 != 5'h0 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_5 | count_6 != 5'h10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_5 | count_6 != 5'h10 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_6 | count_7 != 5'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_6 | count_7 != 5'h0 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_6 | count_7 != 5'h10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_6 | count_7 != 5'h10 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_7 | count_8 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_7 | count_8 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_7 | idle_7 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_7 | idle_7 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_8 | count_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_8 | count_9 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_8 | idle_8 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_8 | idle_8 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_9 | count_10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_9 | count_10 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_9 | idle_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_9 | idle_9 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_10 | count_11 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_10 | count_11 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_10 | idle_10 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_10 | idle_10 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_11 | count_12 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_11 | count_12 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_11 | idle_11 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_11 | idle_11 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_12 | count_13 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_12 | count_13 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_12 | idle_12 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_12 | idle_12 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_13 | count_14 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_13 | count_14 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_13 | idle_13 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_13 | idle_13 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_14 | count_15 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_14 | count_15 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_14 | idle_14 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_14 | idle_14 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_15 | count_16 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_15 | count_16 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_15 | idle_15 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_15 | idle_15 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_16 | count_17 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_16 | count_17 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_16 | idle_16 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_16 | idle_16 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_17 | count_18 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_17 | count_18 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_17 | idle_17 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_17 | idle_17 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_18 | count_19 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_18 | count_19 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_18 | idle_18 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_18 | idle_18 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_19 | count_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_19 | count_20 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_19 | idle_19 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_19 | idle_19 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_20 | count_21 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_20 | count_21 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_20 | idle_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_20 | idle_20 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_21 | count_22 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_21 | count_22 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_21 | idle_21 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_21 | idle_21 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~dec_22 | count_23 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_22 | count_23 | reset)) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~inc_22 | idle_22 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_22 | idle_22 | reset)) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count_7 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  write_6 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  count_6 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  write_5 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  count_5 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  write_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  count_4 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  write_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  count_3 = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  write_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  count_2 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  write_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  count_1 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  write = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  count_23 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  count_22 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  count_21 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  count_20 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  count_19 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  count_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  count_17 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  count_16 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  count_15 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  count_14 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  count_13 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  count_12 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  count_11 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  count_10 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  count_9 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  count_8 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  counter = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  doneAW = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  r_holds_d = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  b_delay = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  r_first = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_denied_r = _RAND_35[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_11(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [12:0] io_in_a_bits_address,
  input  [3:0]  io_in_a_bits_mask,
  input         io_in_a_bits_corrupt,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [2:0]  io_in_c_bits_size,
  input  [6:0]  io_in_c_bits_source,
  input  [12:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [6:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [12:0] _GEN_86 = {{7'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [12:0] _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 13'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_180 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [12:0] _T_183 = io_in_a_bits_address ^ 13'h1000; // @[Parameters.scala 137:31]
  wire [13:0] _T_184 = {1'b0,$signed(_T_183)}; // @[Parameters.scala 137:49]
  wire [13:0] _T_186 = $signed(_T_184) & -14'sh1000; // @[Parameters.scala 137:52]
  wire  _T_187 = $signed(_T_186) == 14'sh0; // @[Parameters.scala 137:67]
  wire  _T_188 = _T_180 & _T_187; // @[Parameters.scala 670:56]
  wire  _T_190 = source_ok & _T_188; // @[Monitor.scala 82:72]
  wire  _T_245 = _source_ok_T_1 & _T_180; // @[Mux.scala 27:72]
  wire  _T_271 = _T_245 & _T_187; // @[Monitor.scala 83:78]
  wire  _T_285 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [3:0] _T_289 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_290 = _T_289 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_294 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18]
  wire  _T_298 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_469 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_482 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_566 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_570 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_578 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_668 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_754 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_755 = io_in_a_bits_mask & _T_754; // @[Monitor.scala 127:31]
  wire  _T_756 = _T_755 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_760 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_842 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_850 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_932 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_940 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1022 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1034 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1038 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1042 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_1046 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_1050 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1054 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1058 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1069 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_1073 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_1086 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1106 = _T_1054 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1115 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1132 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1150 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _source_ok_T_109 = io_in_c_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_115 = io_in_c_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_121 = io_in_c_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_127 = io_in_c_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_133 = io_in_c_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_139 = io_in_c_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_145 = io_in_c_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_151 = io_in_c_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_2 = _source_ok_T_109 | _source_ok_T_115 | _source_ok_T_121 | _source_ok_T_127 | _source_ok_T_133 |
    _source_ok_T_139 | _source_ok_T_145 | _source_ok_T_151; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_7 = 13'h3f << io_in_c_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask_2 = ~_is_aligned_mask_T_7[5:0]; // @[package.scala 234:46]
  wire [12:0] _GEN_87 = {{7'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  wire [12:0] _is_aligned_T_2 = io_in_c_bits_address & _GEN_87; // @[Edges.scala 20:16]
  wire  is_aligned_2 = _is_aligned_T_2 == 13'h0; // @[Edges.scala 20:24]
  wire [12:0] _address_ok_T_5 = io_in_c_bits_address ^ 13'h1000; // @[Parameters.scala 137:31]
  wire [13:0] _address_ok_T_6 = {1'b0,$signed(_address_ok_T_5)}; // @[Parameters.scala 137:49]
  wire [13:0] _address_ok_T_8 = $signed(_address_ok_T_6) & -14'sh1000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_9 = $signed(_address_ok_T_8) == 14'sh0; // @[Parameters.scala 137:67]
  wire  _T_1710 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  wire  _T_1717 = io_in_c_bits_size >= 3'h2; // @[Monitor.scala 245:30]
  wire  _T_1724 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  wire  _T_1732 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  wire  _T_1750 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  wire  _T_1812 = io_in_c_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_1820 = _T_1812 & _address_ok_T_9; // @[Parameters.scala 670:56]
  wire  _T_1822 = source_ok_2 & _T_1820; // @[Monitor.scala 260:78]
  wire  _T_1877 = _source_ok_T_109 & _T_1812; // @[Mux.scala 27:72]
  wire  _T_1903 = _T_1877 & _address_ok_T_9; // @[Monitor.scala 261:78]
  wire  _T_1925 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  wire  _T_2096 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  wire  _T_2106 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  wire  _T_2114 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  wire  _T_2128 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [6:0] source; // @[Monitor.scala 387:22]
  reg [12:0] address; // @[Monitor.scala 388:22]
  wire  _T_2150 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_2151 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_2155 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_2159 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_2163 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_2167 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [6:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_2174 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_2175 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_2179 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_2183 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_2187 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_2195 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  wire  _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  wire [3:0] c_first_beats1_decode = is_aligned_mask_2[5:2]; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  reg [3:0] c_first_counter; // @[Edges.scala 228:27]
  wire [3:0] c_first_counter1 = c_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  c_first = c_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [2:0] size_3; // @[Monitor.scala 514:22]
  reg [6:0] source_3; // @[Monitor.scala 515:22]
  reg [12:0] address_2; // @[Monitor.scala 516:22]
  wire  _T_2226 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  wire  _T_2227 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  wire  _T_2231 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  wire  _T_2235 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  wire  _T_2239 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  wire  _T_2243 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  reg [127:0] inflight; // @[Monitor.scala 611:27]
  reg [511:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [511:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [8:0] _GEN_88 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [9:0] _a_opcode_lookup_T = {{1'd0}, _GEN_88}; // @[Monitor.scala 634:69]
  wire [511:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [511:0] _GEN_89 = {{496'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_89; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[511:1]}; // @[Monitor.scala 634:152]
  wire [511:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [511:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 638:91]
  wire [511:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[511:1]}; // @[Monitor.scala 638:144]
  wire  _T_2249 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [127:0] _a_set_wo_ready_T = 128'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_2252 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [8:0] _GEN_94 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [9:0] _a_opcodes_set_T = {{1'd0}, _GEN_94}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [1026:0] _GEN_95 = {{1023'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [1026:0] _a_opcodes_set_T_1 = _GEN_95 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [1026:0] _GEN_97 = {{1023'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [1026:0] _a_sizes_set_T_1 = _GEN_97 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [127:0] _T_2254 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_2256 = ~_T_2254[0]; // @[Monitor.scala 658:17]
  wire [127:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [1026:0] _GEN_31 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [1026:0] _GEN_32 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_2260 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_2262 = ~_T_1038; // @[Monitor.scala 671:74]
  wire  _T_2263 = io_in_d_valid & d_first_1 & ~_T_1038; // @[Monitor.scala 671:71]
  wire [127:0] _d_clr_wo_ready_T = 128'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1038 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [1038:0] _GEN_99 = {{1023'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [1038:0] _d_opcodes_clr_T_5 = _GEN_99 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [127:0] d_clr = _d_first_T & d_first_1 & _T_2262 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [1038:0] _GEN_35 = _d_first_T & d_first_1 & _T_2262 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_2249 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [127:0] _T_2273 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_2275 = _T_2273[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_2280 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_2281 = io_in_d_bits_opcode == _GEN_44 | _T_2280; // @[Monitor.scala 685:77]
  wire  _T_2285 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_2292 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_2293 = io_in_d_bits_opcode == _GEN_60 | _T_2292; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_102 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_2297 = _GEN_102 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_2307 = _T_2260 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_2262; // @[Monitor.scala 694:116]
  wire  _T_2308 = ~io_in_d_ready; // @[Monitor.scala 695:15]
  wire  _T_2309 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_2316 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [127:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [127:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [127:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [511:0] a_opcodes_set = _GEN_31[511:0];
  wire [511:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [511:0] d_opcodes_clr = _GEN_35[511:0];
  wire [511:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [511:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [511:0] a_sizes_set = _GEN_32[511:0];
  wire [511:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [511:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_2325 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [127:0] inflight_1; // @[Monitor.scala 723:35]
  reg [511:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] c_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] c_first_counter1_1 = c_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  c_first_1 = c_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [511:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [511:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 747:93]
  wire [511:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[511:1]}; // @[Monitor.scala 747:146]
  wire  _T_2335 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  _T_2336 = io_in_c_valid & c_first_1 & _T_2335; // @[Monitor.scala 756:37]
  wire [127:0] _c_set_wo_ready_T = 128'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] c_set_wo_ready = io_in_c_valid & c_first_1 & _T_2335 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 756:71 Monitor.scala 757:22]
  wire  _T_2342 = _c_first_T & c_first_1 & _T_2335; // @[Monitor.scala 760:38]
  wire [3:0] _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  wire [3:0] _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 4'h1; // @[Monitor.scala 763:59]
  wire [8:0] _GEN_109 = {io_in_c_bits_source, 2'h0}; // @[Monitor.scala 764:79]
  wire [9:0] _c_opcodes_set_T = {{1'd0}, _GEN_109}; // @[Monitor.scala 764:79]
  wire [3:0] c_sizes_set_interm = _c_first_T & c_first_1 & _T_2335 ? _c_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 760:72 Monitor.scala 763:28]
  wire [1026:0] _GEN_112 = {{1023'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  wire [1026:0] _c_sizes_set_T_1 = _GEN_112 << _c_opcodes_set_T; // @[Monitor.scala 765:52]
  wire [127:0] _T_2343 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  wire  _T_2345 = ~_T_2343[0]; // @[Monitor.scala 766:17]
  wire [127:0] c_set = _c_first_T & c_first_1 & _T_2335 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 760:72 Monitor.scala 761:28]
  wire [1026:0] _GEN_77 = _c_first_T & c_first_1 & _T_2335 ? _c_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 760:72 Monitor.scala 765:28]
  wire  _T_2349 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  wire  _T_2351 = io_in_d_valid & d_first_2 & _T_1038; // @[Monitor.scala 779:71]
  wire [127:0] d_clr_wo_ready_1 = io_in_d_valid & d_first_2 & _T_1038 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 779:89 Monitor.scala 780:22]
  wire [127:0] d_clr_1 = _d_first_T & d_first_2 & _T_1038 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [1038:0] _GEN_80 = _d_first_T & d_first_2 & _T_1038 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire  _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1 = _T_2336 & io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:88]
  wire [127:0] _T_2359 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire  _T_2361 = _T_2359[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  wire  _T_2365 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_2369 = _GEN_102 == c_size_lookup; // @[Monitor.scala 795:36]
  wire  _T_2378 = _T_2349 & c_first_1 & io_in_c_valid & _same_cycle_resp_T_8 & _T_1038; // @[Monitor.scala 799:116]
  wire  _T_2380 = _T_2308 | io_in_c_ready; // @[Monitor.scala 800:32]
  wire  _T_2384 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  wire  _T_2385 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  wire [127:0] _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  wire [127:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [127:0] _inflight_T_5 = _inflight_T_3 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [511:0] d_opcodes_clr_1 = _GEN_80[511:0];
  wire [511:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [511:0] c_sizes_set = _GEN_77[511:0];
  wire [511:0] _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  wire [511:0] _inflight_sizes_T_5 = _inflight_sizes_T_3 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_2394 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [3:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_3 = d_first_counter_3 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 4'h0; // @[Edges.scala 230:25]
  wire  _T_2406 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_2407 = _d_first_T & d_first_3 & _T_2406; // @[Monitor.scala 829:38]
  wire  _T_2410 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = _d_first_T & d_first_3 & _T_2406 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  d_set = _GEN_84[0];
  wire  _T_2417 = d_set | inflight_2; // @[Monitor.scala 837:24]
  wire [1:0] _GEN_85 = io_in_e_valid ? 2'h1 : 2'h0; // @[Monitor.scala 835:73 Monitor.scala 836:13]
  wire  e_clr = _GEN_85[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 4'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      opcode_3 <= io_in_c_bits_opcode; // @[Monitor.scala 525:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      param_3 <= io_in_c_bits_param; // @[Monitor.scala 526:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      size_3 <= io_in_c_bits_size; // @[Monitor.scala 527:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      source_3 <= io_in_c_bits_source; // @[Monitor.scala 528:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      address_2 <= io_in_c_bits_address; // @[Monitor.scala 529:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 128'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 512'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 512'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 128'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 512'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first_1) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 4'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_c_first_T | _d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= (inflight_2 | d_set) & ~e_clr; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 4'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_271 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_271 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_285 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_285 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_290 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_290 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_294 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_294 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_271 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_271 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_285 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_285 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_469 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_469 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_290 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_290 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_294 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_294 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_188 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_188 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_566 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_566 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_294 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_294 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_566 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_566 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_566 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_566 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_756 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_756 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_842 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_842 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_932 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_932 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_1022 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_1022 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_294 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_294 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1034 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1034 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1042 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1042 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1046 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1046 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1054 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1054 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1042 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1042 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1069 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1069 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1073 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1073 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1042 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1042 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1069 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1069 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1073 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1073 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1106 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(_T_1046 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(_T_1046 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(_T_1050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(_T_1050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(_T_1046 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(_T_1046 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(_T_1106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(_T_1106 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(_T_1046 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(_T_1046 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(_T_1050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(_T_1050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_T_1717 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_T_1717 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_T_1724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_T_1724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_T_1717 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_T_1717 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_T_1724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_T_1724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1822 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1822 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1903 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1903 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1717 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1717 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid report param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1822 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1822 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1903 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1903 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1717 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1717 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(_T_2106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(_T_2106 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(_T_2106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(_T_2106 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(_T_2106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(_T_2106 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2151 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2151 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2155 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2155 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2159 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2159 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2163 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2163 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2167 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2167 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2175 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2175 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2179 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2179 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2183 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2183 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2187 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2187 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2195 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2195 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2227 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2227 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2235 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2235 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2239 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2239 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2243 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2243 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2252 & ~(_T_2256 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2252 & ~(_T_2256 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & ~(_T_2275 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & ~(_T_2275 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & same_cycle_resp & ~(_T_2281 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & same_cycle_resp & ~(_T_2281 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & same_cycle_resp & ~(_T_2285 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & same_cycle_resp & ~(_T_2285 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & ~same_cycle_resp & ~(_T_2293 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & ~same_cycle_resp & ~(_T_2293 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & ~same_cycle_resp & ~(_T_2297 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & ~same_cycle_resp & ~(_T_2297 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2307 & ~(_T_2309 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2307 & ~(_T_2309 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2316 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2316 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2325 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2325 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2342 & ~(_T_2345 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel re-used a source ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2342 & ~(_T_2345 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2351 & ~(_T_2361 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2351 & ~(_T_2361 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2351 & same_cycle_resp_1 & ~(_T_2365 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2351 & same_cycle_resp_1 & ~(_T_2365 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2351 & ~same_cycle_resp_1 & ~(_T_2369 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2351 & ~same_cycle_resp_1 & ~(_T_2369 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2378 & ~(_T_2380 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2378 & ~(_T_2380 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2384 & ~(_T_2385 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2384 & ~(_T_2385 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2394 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2394 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2407 & ~(_T_2410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2407 & ~(_T_2410 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & ~(_T_2417 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:154:12)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & ~(_T_2417 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  c_first_counter = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  opcode_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  param_3 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  size_3 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  source_3 = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  address_2 = _RAND_17[12:0];
  _RAND_18 = {4{`RANDOM}};
  inflight = _RAND_18[127:0];
  _RAND_19 = {16{`RANDOM}};
  inflight_opcodes = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  inflight_sizes = _RAND_20[511:0];
  _RAND_21 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  watchdog = _RAND_23[31:0];
  _RAND_24 = {4{`RANDOM}};
  inflight_1 = _RAND_24[127:0];
  _RAND_25 = {16{`RANDOM}};
  inflight_sizes_1 = _RAND_25[511:0];
  _RAND_26 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  watchdog_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inflight_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_30[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_18(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [2:0] io_enq_bits_size,
  input  [6:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_size,
  output [6:0] io_deq_bits_source
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_source [0:0]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign ram_opcode_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = 1'h0;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = 1'h0;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[6:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_19(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [2:0] io_enq_bits_param,
  input  [2:0] io_enq_bits_size,
  input  [6:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [2:0] io_deq_bits_size,
  output [6:0] io_deq_bits_source
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_param [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_source [0:0]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 224:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign ram_opcode_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = 1'h0;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = 1'h0;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = 1'h0;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[6:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLError_2(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [12:0] auto_in_a_bits_address,
  input  [3:0]  auto_in_a_bits_mask,
  input         auto_in_a_bits_corrupt,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [2:0]  auto_in_c_bits_size,
  input  [6:0]  auto_in_c_bits_source,
  input  [12:0] auto_in_c_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output        auto_in_d_bits_corrupt,
  input         auto_in_e_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [12:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [12:0] monitor_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_valid; // @[Nodes.scala 24:25]
  wire  a_clock; // @[Decoupled.scala 296:21]
  wire  a_reset; // @[Decoupled.scala 296:21]
  wire  a_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  a_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] a_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] a_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [6:0] a_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire  a_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  a_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] a_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] a_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [6:0] a_io_deq_bits_source; // @[Decoupled.scala 296:21]
  wire  c_clock; // @[Decoupled.scala 296:21]
  wire  c_reset; // @[Decoupled.scala 296:21]
  wire  c_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  c_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] c_io_enq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] c_io_enq_bits_param; // @[Decoupled.scala 296:21]
  wire [2:0] c_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire [6:0] c_io_enq_bits_source; // @[Decoupled.scala 296:21]
  wire  c_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  c_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [2:0] c_io_deq_bits_opcode; // @[Decoupled.scala 296:21]
  wire [2:0] c_io_deq_bits_param; // @[Decoupled.scala 296:21]
  wire [2:0] c_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire [6:0] c_io_deq_bits_source; // @[Decoupled.scala 296:21]
  reg  idle; // @[Error.scala 44:23]
  wire  _a_last_T = a_io_deq_ready & a_io_deq_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _a_last_beats1_decode_T_1 = 13'h3f << a_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] _a_last_beats1_decode_T_3 = ~_a_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] a_last_beats1_decode = _a_last_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  a_last_beats1_opdata = ~a_io_deq_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [3:0] a_last_beats1 = a_last_beats1_opdata ? a_last_beats1_decode : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] a_last_counter; // @[Edges.scala 228:27]
  wire [3:0] a_last_counter1 = a_last_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_last_first = a_last_counter == 4'h0; // @[Edges.scala 230:25]
  wire  a_last = a_last_counter == 4'h1 | a_last_beats1 == 4'h0; // @[Edges.scala 231:37]
  reg [3:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle_1 = beatsLeft == 4'h0; // @[Arbiter.scala 88:28]
  wire  da_valid = a_io_deq_valid & a_last & idle; // @[Error.scala 51:35]
  reg [3:0] c_last_counter; // @[Edges.scala 228:27]
  wire  c_last_beats1_opdata = c_io_deq_bits_opcode[0]; // @[Edges.scala 101:36]
  wire [12:0] _c_last_beats1_decode_T_1 = 13'h3f << c_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] _c_last_beats1_decode_T_3 = ~_c_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] c_last_beats1_decode = _c_last_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire [3:0] c_last_beats1 = c_last_beats1_opdata ? c_last_beats1_decode : 4'h0; // @[Edges.scala 220:14]
  wire  c_last = c_last_counter == 4'h1 | c_last_beats1 == 4'h0; // @[Edges.scala 231:37]
  wire  dc_valid = c_io_deq_valid & c_last; // @[Error.scala 74:27]
  wire [1:0] _readys_T = {da_valid,dc_valid}; // @[Cat.scala 30:58]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[package.scala 244:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[Arbiter.scala 16:61]
  wire  readys_1 = _readys_T_7[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle_1 ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_in_d_ready & allowed_1; // @[Arbiter.scala 123:31]
  wire  _T = out_1_ready & da_valid; // @[Decoupled.scala 40:37]
  wire [2:0] da_bits_size = a_io_deq_bits_size; // @[Error.scala 43:18 Error.scala 55:21]
  wire [12:0] _beats1_decode_T_1 = 13'h3f << da_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] beats1_decode = _beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire [2:0] _GEN_4 = 3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_5 = 3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_4; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_6 = 3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_5; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_7 = 3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_6; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] _GEN_8 = 3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_7; // @[Error.scala 53:21 Error.scala 53:21]
  wire [2:0] da_bits_opcode = 3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8; // @[Error.scala 53:21 Error.scala 53:21]
  wire  beats1_opdata = da_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [3:0] beats1 = beats1_opdata ? beats1_decode : 4'h0; // @[Edges.scala 220:14]
  reg [3:0] counter; // @[Edges.scala 228:27]
  wire [3:0] counter1 = counter - 4'h1; // @[Edges.scala 229:28]
  wire  da_first = counter == 4'h0; // @[Edges.scala 230:25]
  wire  da_last = counter == 4'h1 | beats1 == 4'h0; // @[Edges.scala 231:37]
  wire  _c_last_T = c_io_deq_ready & c_io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] c_last_counter1 = c_last_counter - 4'h1; // @[Edges.scala 229:28]
  wire  c_last_first = c_last_counter == 4'h0; // @[Edges.scala 230:25]
  wire  readys_0 = _readys_T_7[0]; // @[Arbiter.scala 95:86]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  allowed_0 = idle_1 ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  out_ready = auto_in_d_ready & allowed_0; // @[Arbiter.scala 123:31]
  wire [2:0] dc_bits_size = c_io_deq_bits_size; // @[Error.scala 64:20 Error.scala 79:23]
  wire  _GEN_12 = _T & da_bits_opcode == 3'h4 ? 1'h0 : idle; // @[Error.scala 70:52 Error.scala 70:59 Error.scala 44:23]
  wire  _GEN_13 = auto_in_e_valid | _GEN_12; // @[Error.scala 71:26 Error.scala 71:33]
  wire [1:0] _GEN_15 = 2'h1 == c_io_deq_bits_param[1:0] ? 2'h2 : 2'h1; // @[Error.scala 78:23 Error.scala 78:23]
  wire [1:0] dc_bits_param = 2'h2 == c_io_deq_bits_param[1:0] ? 2'h2 : _GEN_15; // @[Error.scala 78:23 Error.scala 78:23]
  wire  latch = idle_1 & auto_in_d_ready; // @[Arbiter.scala 89:24]
  wire  earlyWinner_0 = readys_0 & dc_valid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1 = readys_1 & da_valid; // @[Arbiter.scala 97:79]
  wire  _prefixOR_T = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 104:53]
  wire  _T_21 = dc_valid | da_valid; // @[Arbiter.scala 107:36]
  wire  _T_22 = ~(dc_valid | da_valid); // @[Arbiter.scala 107:15]
  wire  muxStateEarly_0 = idle_1 ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly_1 = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & dc_valid | state_1 & da_valid; // @[Mux.scala 27:72]
  wire  sink_ACancel_earlyValid = idle_1 ? _T_21 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 50:33]
  wire [3:0] _GEN_17 = {{3'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [3:0] _beatsLeft_T_4 = beatsLeft - _GEN_17; // @[Arbiter.scala 113:52]
  wire [6:0] dc_bits_source = c_io_deq_bits_source; // @[Error.scala 64:20 Error.scala 80:23]
  wire [6:0] _T_47 = muxStateEarly_0 ? dc_bits_source : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] da_bits_source = a_io_deq_bits_source; // @[Error.scala 43:18 Error.scala 56:21]
  wire [6:0] _T_48 = muxStateEarly_1 ? da_bits_source : 7'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_50 = muxStateEarly_0 ? dc_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_51 = muxStateEarly_1 ? da_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_56 = muxStateEarly_0 ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_57 = muxStateEarly_1 ? da_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  TLMonitor_11 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_c_ready(monitor_io_in_c_ready),
    .io_in_c_valid(monitor_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_io_in_c_bits_address),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),
    .io_in_e_valid(monitor_io_in_e_valid)
  );
  Queue_18 a ( // @[Decoupled.scala 296:21]
    .clock(a_clock),
    .reset(a_reset),
    .io_enq_ready(a_io_enq_ready),
    .io_enq_valid(a_io_enq_valid),
    .io_enq_bits_opcode(a_io_enq_bits_opcode),
    .io_enq_bits_size(a_io_enq_bits_size),
    .io_enq_bits_source(a_io_enq_bits_source),
    .io_deq_ready(a_io_deq_ready),
    .io_deq_valid(a_io_deq_valid),
    .io_deq_bits_opcode(a_io_deq_bits_opcode),
    .io_deq_bits_size(a_io_deq_bits_size),
    .io_deq_bits_source(a_io_deq_bits_source)
  );
  Queue_19 c ( // @[Decoupled.scala 296:21]
    .clock(c_clock),
    .reset(c_reset),
    .io_enq_ready(c_io_enq_ready),
    .io_enq_valid(c_io_enq_valid),
    .io_enq_bits_opcode(c_io_enq_bits_opcode),
    .io_enq_bits_param(c_io_enq_bits_param),
    .io_enq_bits_size(c_io_enq_bits_size),
    .io_enq_bits_source(c_io_enq_bits_source),
    .io_deq_ready(c_io_deq_ready),
    .io_deq_valid(c_io_deq_valid),
    .io_deq_bits_opcode(c_io_deq_bits_opcode),
    .io_deq_bits_param(c_io_deq_bits_param),
    .io_deq_bits_size(c_io_deq_bits_size),
    .io_deq_bits_source(c_io_deq_bits_source)
  );
  assign auto_in_a_ready = a_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign auto_in_c_ready = c_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign auto_in_d_valid = idle_1 ? _T_21 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_in_d_bits_opcode = _T_56 | _T_57; // @[Mux.scala 27:72]
  assign auto_in_d_bits_param = muxStateEarly_0 ? dc_bits_param : 2'h0; // @[Mux.scala 27:72]
  assign auto_in_d_bits_size = _T_50 | _T_51; // @[Mux.scala 27:72]
  assign auto_in_d_bits_source = _T_47 | _T_48; // @[Mux.scala 27:72]
  assign auto_in_d_bits_denied = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  assign auto_in_d_bits_corrupt = muxStateEarly_1 & beats1_opdata; // @[Mux.scala 27:72]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = a_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_ready = c_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 299:17]
  assign monitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = idle_1 ? _T_21 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign monitor_io_in_d_bits_opcode = _T_56 | _T_57; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_param = muxStateEarly_0 ? dc_bits_param : 2'h0; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_size = _T_50 | _T_51; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_source = _T_47 | _T_48; // @[Mux.scala 27:72]
  assign monitor_io_in_d_bits_denied = idle_1 ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  assign monitor_io_in_d_bits_corrupt = muxStateEarly_1 & beats1_opdata; // @[Mux.scala 27:72]
  assign monitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_clock = clock;
  assign a_reset = reset;
  assign a_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_deq_ready = out_1_ready & da_last & idle | ~a_last; // @[Error.scala 50:46]
  assign c_clock = clock;
  assign c_reset = reset;
  assign c_io_enq_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign c_io_enq_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign c_io_enq_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign c_io_enq_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign c_io_enq_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign c_io_deq_ready = out_ready | ~c_last; // @[Error.scala 73:40]
  always @(posedge clock) begin
    idle <= reset | _GEN_13; // @[Error.scala 44:23 Error.scala 44:23]
    if (reset) begin // @[Edges.scala 228:27]
      a_last_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_last_T) begin // @[Edges.scala 234:17]
      if (a_last_first) begin // @[Edges.scala 235:21]
        if (a_last_beats1_opdata) begin // @[Edges.scala 220:14]
          a_last_counter <= a_last_beats1_decode;
        end else begin
          a_last_counter <= 4'h0;
        end
      end else begin
        a_last_counter <= a_last_counter1;
      end
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 4'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin // @[Arbiter.scala 113:23]
      if (earlyWinner_1) begin // @[Arbiter.scala 111:73]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          beatsLeft <= beats1_decode;
        end else begin
          beatsLeft <= 4'h0;
        end
      end else begin
        beatsLeft <= 4'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_last_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_c_last_T) begin // @[Edges.scala 234:17]
      if (c_last_first) begin // @[Edges.scala 235:21]
        if (c_last_beats1_opdata) begin // @[Edges.scala 220:14]
          c_last_counter <= c_last_beats1_decode;
        end else begin
          c_last_counter <= 4'h0;
        end
      end else begin
        c_last_counter <= c_last_counter1;
      end
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin // @[Arbiter.scala 117:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_T) begin // @[Edges.scala 234:17]
      if (da_first) begin // @[Edges.scala 235:21]
        if (beats1_opdata) begin // @[Edges.scala 220:14]
          counter <= beats1_decode;
        end else begin
          counter <= 4'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin // @[Arbiter.scala 117:30]
      state_0 <= earlyWinner_0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(idle | da_first | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Error.scala:49 assert (idle || da_first) // we only send Grant, never GrantData => simplified flow control below\n"
            ); // @[Error.scala 49:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(idle | da_first | reset)) begin
          $fatal; // @[Error.scala 49:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(dc_valid | da_valid) | _prefixOR_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(dc_valid | da_valid) | _prefixOR_T | reset)) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_22 | _T_21 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_22 | _T_21 | reset)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  idle = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  a_last_counter = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  beatsLeft = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  c_last_counter = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  state_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  counter = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  state_0 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_12(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [2:0]  io_in_c_bits_size,
  input  [6:0]  io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [6:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input         io_in_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_86 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_2 = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_3 = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_4 = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_5 = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_lo = mask_acc_2 | mask_size_2 & mask_eq_6; // @[Misc.scala 214:29]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_hi = mask_acc_2 | mask_size_2 & mask_eq_7; // @[Misc.scala 214:29]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_lo = mask_acc_3 | mask_size_2 & mask_eq_8; // @[Misc.scala 214:29]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_hi = mask_acc_3 | mask_size_2 & mask_eq_9; // @[Misc.scala 214:29]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_lo = mask_acc_4 | mask_size_2 & mask_eq_10; // @[Misc.scala 214:29]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_hi = mask_acc_4 | mask_size_2 & mask_eq_11; // @[Misc.scala 214:29]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_lo = mask_acc_5 | mask_size_2 & mask_eq_12; // @[Misc.scala 214:29]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_hi = mask_acc_5 | mask_size_2 & mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire [31:0] _T_180 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_181 = {1'b0,$signed(_T_180)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_183 = $signed(_T_181) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_184 = $signed(_T_183) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_185 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_186 = {1'b0,$signed(_T_185)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_188 = $signed(_T_186) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_189 = $signed(_T_188) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_190 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_191 = {1'b0,$signed(_T_190)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_193 = $signed(_T_191) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_194 = $signed(_T_193) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_195 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_196 = {1'b0,$signed(_T_195)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_198 = $signed(_T_196) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_199 = $signed(_T_198) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_200 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_201 = {1'b0,$signed(_T_200)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_203 = $signed(_T_201) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_204 = $signed(_T_203) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_211 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_214 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_215 = {1'b0,$signed(_T_214)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_217 = $signed(_T_215) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_218 = $signed(_T_217) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_219 = _T_211 & _T_218; // @[Parameters.scala 670:56]
  wire  _T_222 = source_ok & _T_219; // @[Monitor.scala 82:72]
  wire  _T_277 = _source_ok_T_1 & _T_211; // @[Mux.scala 27:72]
  wire  _T_330 = _T_218 | _T_184 | _T_189 | _T_194 | _T_199 | _T_204; // @[Parameters.scala 671:42]
  wire  _T_333 = _T_277 & _T_330; // @[Monitor.scala 83:78]
  wire  _T_347 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [7:0] _T_351 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_352 = _T_351 == 8'h0; // @[Monitor.scala 88:31]
  wire  _T_360 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_593 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_606 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_709 = _T_211 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_720 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_724 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_732 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_834 = source_ok & _T_709; // @[Monitor.scala 115:71]
  wire  _T_852 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [7:0] _T_968 = ~mask; // @[Monitor.scala 127:33]
  wire [7:0] _T_969 = io_in_a_bits_mask & _T_968; // @[Monitor.scala 127:31]
  wire  _T_970 = _T_969 == 8'h0; // @[Monitor.scala 127:40]
  wire  _T_974 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_1036 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_1074 = _T_1036 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_1076 = source_ok & _T_1074; // @[Monitor.scala 131:74]
  wire  _T_1086 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_1094 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_1206 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_1214 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1328 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1340 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1344 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1348 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27]
  wire  _T_1352 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_1356 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1360 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1364 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1375 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_1379 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_1392 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1412 = _T_1360 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1421 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1438 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1456 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _source_ok_T_109 = io_in_c_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_115 = io_in_c_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_121 = io_in_c_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_127 = io_in_c_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_133 = io_in_c_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_139 = io_in_c_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_145 = io_in_c_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_151 = io_in_c_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_2 = _source_ok_T_109 | _source_ok_T_115 | _source_ok_T_121 | _source_ok_T_127 | _source_ok_T_133 |
    _source_ok_T_139 | _source_ok_T_145 | _source_ok_T_151; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_7 = 13'h3f << io_in_c_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask_2 = ~_is_aligned_mask_T_7[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_87 = {{26'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T_2 = io_in_c_bits_address & _GEN_87; // @[Edges.scala 20:16]
  wire  is_aligned_2 = _is_aligned_T_2 == 32'h0; // @[Edges.scala 20:24]
  wire [31:0] _address_ok_T_34 = io_in_c_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_35 = {1'b0,$signed(_address_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_37 = $signed(_address_ok_T_35) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_38 = $signed(_address_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_39 = io_in_c_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_40 = {1'b0,$signed(_address_ok_T_39)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_42 = $signed(_address_ok_T_40) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_43 = $signed(_address_ok_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_44 = io_in_c_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_45 = {1'b0,$signed(_address_ok_T_44)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_47 = $signed(_address_ok_T_45) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_48 = $signed(_address_ok_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_49 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_50 = {1'b0,$signed(_address_ok_T_49)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_52 = $signed(_address_ok_T_50) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_53 = $signed(_address_ok_T_52) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_54 = io_in_c_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_55 = {1'b0,$signed(_address_ok_T_54)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_57 = $signed(_address_ok_T_55) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_58 = $signed(_address_ok_T_57) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _address_ok_T_62 = _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 | _address_ok_T_58; // @[Parameters.scala 598:92]
  wire [31:0] _address_ok_T_63 = io_in_c_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_64 = {1'b0,$signed(_address_ok_T_63)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_66 = $signed(_address_ok_T_64) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_67 = $signed(_address_ok_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  wire  address_ok_1 = _address_ok_T_62 | _address_ok_T_67; // @[Parameters.scala 622:64]
  wire  _T_2226 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  wire  _T_2233 = io_in_c_bits_size >= 3'h3; // @[Monitor.scala 245:30]
  wire  _T_2240 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  wire  _T_2248 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  wire  _T_2266 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  wire  _T_2359 = io_in_c_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_2367 = _T_2359 & _address_ok_T_67; // @[Parameters.scala 670:56]
  wire  _T_2370 = source_ok_2 & _T_2367; // @[Monitor.scala 260:78]
  wire  _T_2425 = _source_ok_T_109 & _T_2359; // @[Mux.scala 27:72]
  wire  _T_2478 = _address_ok_T_67 | _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 |
    _address_ok_T_58; // @[Parameters.scala 671:42]
  wire  _T_2481 = _T_2425 & _T_2478; // @[Monitor.scala 261:78]
  wire  _T_2503 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  wire  _T_2736 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  wire  _T_2746 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  wire  _T_2754 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  wire  _T_2768 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  wire  sink_ok_1 = io_in_e_bits_sink < 1'h1; // @[Monitor.scala 364:31]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [6:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_2790 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_2791 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_2795 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_2799 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_2803 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_2807 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [6:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_2814 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_2815 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_2819 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_2823 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_2827 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_2835 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  wire  _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  wire [2:0] c_first_beats1_decode = is_aligned_mask_2[5:3]; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  reg [2:0] c_first_counter; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1 = c_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  c_first = c_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [2:0] size_3; // @[Monitor.scala 514:22]
  reg [6:0] source_3; // @[Monitor.scala 515:22]
  reg [31:0] address_2; // @[Monitor.scala 516:22]
  wire  _T_2866 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  wire  _T_2867 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  wire  _T_2871 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  wire  _T_2875 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  wire  _T_2879 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  wire  _T_2883 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  reg [127:0] inflight; // @[Monitor.scala 611:27]
  reg [511:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [511:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  wire [8:0] _GEN_88 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [9:0] _a_opcode_lookup_T = {{1'd0}, _GEN_88}; // @[Monitor.scala 634:69]
  wire [511:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [511:0] _GEN_89 = {{496'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_89; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[511:1]}; // @[Monitor.scala 634:152]
  wire [511:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [511:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 638:91]
  wire [511:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[511:1]}; // @[Monitor.scala 638:144]
  wire  _T_2889 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [127:0] _a_set_wo_ready_T = 128'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_2892 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [8:0] _GEN_94 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [9:0] _a_opcodes_set_T = {{1'd0}, _GEN_94}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [1026:0] _GEN_95 = {{1023'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [1026:0] _a_opcodes_set_T_1 = _GEN_95 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [1026:0] _GEN_97 = {{1023'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [1026:0] _a_sizes_set_T_1 = _GEN_97 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [127:0] _T_2894 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_2896 = ~_T_2894[0]; // @[Monitor.scala 658:17]
  wire [127:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [1026:0] _GEN_31 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [1026:0] _GEN_32 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_2900 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_2902 = ~_T_1344; // @[Monitor.scala 671:74]
  wire  _T_2903 = io_in_d_valid & d_first_1 & ~_T_1344; // @[Monitor.scala 671:71]
  wire [127:0] _d_clr_wo_ready_T = 128'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1344 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [1038:0] _GEN_99 = {{1023'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [1038:0] _d_opcodes_clr_T_5 = _GEN_99 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [127:0] d_clr = _d_first_T & d_first_1 & _T_2902 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [1038:0] _GEN_35 = _d_first_T & d_first_1 & _T_2902 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_2889 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [127:0] _T_2913 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_2915 = _T_2913[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_2920 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_2921 = io_in_d_bits_opcode == _GEN_44 | _T_2920; // @[Monitor.scala 685:77]
  wire  _T_2925 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_2932 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_2933 = io_in_d_bits_opcode == _GEN_60 | _T_2932; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_102 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_2937 = _GEN_102 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_2947 = _T_2900 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_2902; // @[Monitor.scala 694:116]
  wire  _T_2948 = ~io_in_d_ready; // @[Monitor.scala 695:15]
  wire  _T_2949 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_2956 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [127:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [127:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [127:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [511:0] a_opcodes_set = _GEN_31[511:0];
  wire [511:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [511:0] d_opcodes_clr = _GEN_35[511:0];
  wire [511:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [511:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [511:0] a_sizes_set = _GEN_32[511:0];
  wire [511:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [511:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_2965 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [127:0] inflight_1; // @[Monitor.scala 723:35]
  reg [511:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [2:0] c_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1_1 = c_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  c_first_1 = c_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25]
  wire [511:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [511:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 747:93]
  wire [511:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[511:1]}; // @[Monitor.scala 747:146]
  wire  _T_2975 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  _T_2976 = io_in_c_valid & c_first_1 & _T_2975; // @[Monitor.scala 756:37]
  wire [127:0] _c_set_wo_ready_T = 128'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] c_set_wo_ready = io_in_c_valid & c_first_1 & _T_2975 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 756:71 Monitor.scala 757:22]
  wire  _T_2982 = _c_first_T & c_first_1 & _T_2975; // @[Monitor.scala 760:38]
  wire [3:0] _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  wire [3:0] _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 4'h1; // @[Monitor.scala 763:59]
  wire [8:0] _GEN_109 = {io_in_c_bits_source, 2'h0}; // @[Monitor.scala 764:79]
  wire [9:0] _c_opcodes_set_T = {{1'd0}, _GEN_109}; // @[Monitor.scala 764:79]
  wire [3:0] c_sizes_set_interm = _c_first_T & c_first_1 & _T_2975 ? _c_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 760:72 Monitor.scala 763:28]
  wire [1026:0] _GEN_112 = {{1023'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  wire [1026:0] _c_sizes_set_T_1 = _GEN_112 << _c_opcodes_set_T; // @[Monitor.scala 765:52]
  wire [127:0] _T_2983 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  wire  _T_2985 = ~_T_2983[0]; // @[Monitor.scala 766:17]
  wire [127:0] c_set = _c_first_T & c_first_1 & _T_2975 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 760:72 Monitor.scala 761:28]
  wire [1026:0] _GEN_77 = _c_first_T & c_first_1 & _T_2975 ? _c_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 760:72 Monitor.scala 765:28]
  wire  _T_2989 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  wire  _T_2991 = io_in_d_valid & d_first_2 & _T_1344; // @[Monitor.scala 779:71]
  wire [127:0] d_clr_wo_ready_1 = io_in_d_valid & d_first_2 & _T_1344 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 779:89 Monitor.scala 780:22]
  wire [127:0] d_clr_1 = _d_first_T & d_first_2 & _T_1344 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [1038:0] _GEN_80 = _d_first_T & d_first_2 & _T_1344 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire  _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1 = _T_2976 & io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:88]
  wire [127:0] _T_2999 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire  _T_3001 = _T_2999[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  wire  _T_3005 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_3009 = _GEN_102 == c_size_lookup; // @[Monitor.scala 795:36]
  wire  _T_3018 = _T_2989 & c_first_1 & io_in_c_valid & _same_cycle_resp_T_8 & _T_1344; // @[Monitor.scala 799:116]
  wire  _T_3020 = _T_2948 | io_in_c_ready; // @[Monitor.scala 800:32]
  wire  _T_3024 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  wire  _T_3025 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  wire [127:0] _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  wire [127:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [127:0] _inflight_T_5 = _inflight_T_3 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [511:0] d_opcodes_clr_1 = _GEN_80[511:0];
  wire [511:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [511:0] c_sizes_set = _GEN_77[511:0];
  wire [511:0] _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  wire [511:0] _inflight_sizes_T_5 = _inflight_sizes_T_3 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_3034 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [2:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_3 = d_first_counter_3 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 3'h0; // @[Edges.scala 230:25]
  wire  _T_3046 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_3047 = _d_first_T & d_first_3 & _T_3046; // @[Monitor.scala 829:38]
  wire  _T_3050 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = _d_first_T & d_first_3 & _T_3046 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  _T_3054 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _e_clr_T = 2'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  wire  d_set = _GEN_84[0];
  wire  _T_3058 = (d_set | inflight_2) >> io_in_e_bits_sink; // @[Monitor.scala 837:35]
  wire [1:0] _GEN_85 = _T_3054 ? _e_clr_T : 2'h0; // @[Monitor.scala 835:73 Monitor.scala 836:13]
  wire  e_clr = _GEN_85[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 3'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      opcode_3 <= io_in_c_bits_opcode; // @[Monitor.scala 525:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      param_3 <= io_in_c_bits_param; // @[Monitor.scala 526:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      size_3 <= io_in_c_bits_size; // @[Monitor.scala 527:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      source_3 <= io_in_c_bits_source; // @[Monitor.scala 528:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      address_2 <= io_in_c_bits_address; // @[Monitor.scala 529:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 128'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 512'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 512'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 128'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 512'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first_1) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 3'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_c_first_T | _d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= (inflight_2 | d_set) & ~e_clr; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 3'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1328 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1328 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1340 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1340 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1348 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1348 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1360 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1360 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1348 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1348 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1375 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1375 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1379 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1379 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1348 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1348 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1375 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1375 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1379 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1379 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1412 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1412 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(_T_1412 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(_T_1412 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(_T_2233 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(_T_2233 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(_T_2240 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(_T_2240 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(_T_2233 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(_T_2233 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(_T_2240 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(_T_2240 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2370 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2370 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2481 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2481 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2233 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2233 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2240 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid report param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2240 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2370 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2370 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2481 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2481 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2233 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2233 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2240 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2240 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(_T_2746 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(_T_2746 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(_T_2746 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(_T_2746 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(_T_2746 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(_T_2746 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channels carries invalid sink ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2791 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2791 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2795 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2795 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2799 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2799 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2803 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2803 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2807 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2807 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2815 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2815 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2819 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2819 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2823 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2823 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2827 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2827 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2835 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2835 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2867 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2867 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2871 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2871 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2875 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2875 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2879 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2879 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2883 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2883 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2892 & ~(_T_2896 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2892 & ~(_T_2896 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & ~(_T_2915 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & ~(_T_2915 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & same_cycle_resp & ~(_T_2921 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & same_cycle_resp & ~(_T_2921 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & same_cycle_resp & ~(_T_2925 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & same_cycle_resp & ~(_T_2925 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & ~same_cycle_resp & ~(_T_2933 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & ~same_cycle_resp & ~(_T_2933 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & ~same_cycle_resp & ~(_T_2937 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & ~same_cycle_resp & ~(_T_2937 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2947 & ~(_T_2949 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2947 & ~(_T_2949 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2956 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2956 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2965 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2965 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2982 & ~(_T_2985 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel re-used a source ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2982 & ~(_T_2985 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2991 & ~(_T_3001 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2991 & ~(_T_3001 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2991 & same_cycle_resp_1 & ~(_T_3005 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2991 & same_cycle_resp_1 & ~(_T_3005 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2991 & ~same_cycle_resp_1 & ~(_T_3009 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2991 & ~same_cycle_resp_1 & ~(_T_3009 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3018 & ~(_T_3020 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3018 & ~(_T_3020 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3024 & ~(_T_3025 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3024 & ~(_T_3025 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_3034 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_3034 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3047 & ~(_T_3050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3047 & ~(_T_3050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3054 & ~(_T_3058 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:47)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3054 & ~(_T_3058 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  c_first_counter = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  opcode_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  param_3 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  size_3 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  source_3 = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  address_2 = _RAND_17[31:0];
  _RAND_18 = {4{`RANDOM}};
  inflight = _RAND_18[127:0];
  _RAND_19 = {16{`RANDOM}};
  inflight_opcodes = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  inflight_sizes = _RAND_20[511:0];
  _RAND_21 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  watchdog = _RAND_23[31:0];
  _RAND_24 = {4{`RANDOM}};
  inflight_1 = _RAND_24[127:0];
  _RAND_25 = {16{`RANDOM}};
  inflight_sizes_1 = _RAND_25[511:0];
  _RAND_26 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  watchdog_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inflight_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_30[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLAtomicAutomata(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [2:0]  auto_in_c_bits_size,
  input  [6:0]  auto_in_c_bits_source,
  input  [31:0] auto_in_c_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  output        auto_in_e_ready,
  input         auto_in_e_valid,
  input         auto_in_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [2:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_a_bits_corrupt,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [2:0]  auto_out_c_bits_size,
  output [6:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [2:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output        auto_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_bits_sink; // @[Nodes.scala 24:25]
  reg [1:0] cam_s_0_state; // @[AtomicAutomata.scala 76:28]
  reg [2:0] cam_a_0_bits_opcode; // @[AtomicAutomata.scala 77:24]
  reg [2:0] cam_a_0_bits_param; // @[AtomicAutomata.scala 77:24]
  reg [2:0] cam_a_0_bits_size; // @[AtomicAutomata.scala 77:24]
  reg [6:0] cam_a_0_bits_source; // @[AtomicAutomata.scala 77:24]
  reg [31:0] cam_a_0_bits_address; // @[AtomicAutomata.scala 77:24]
  reg [7:0] cam_a_0_bits_mask; // @[AtomicAutomata.scala 77:24]
  reg [63:0] cam_a_0_bits_data; // @[AtomicAutomata.scala 77:24]
  reg  cam_a_0_fifoId; // @[AtomicAutomata.scala 77:24]
  reg [3:0] cam_a_0_lut; // @[AtomicAutomata.scala 77:24]
  reg [63:0] cam_d_0_data; // @[AtomicAutomata.scala 78:24]
  reg  cam_d_0_denied; // @[AtomicAutomata.scala 78:24]
  reg  cam_d_0_corrupt; // @[AtomicAutomata.scala 78:24]
  wire  cam_free_0 = cam_s_0_state == 2'h0; // @[AtomicAutomata.scala 80:44]
  wire  cam_amo_0 = cam_s_0_state == 2'h2; // @[AtomicAutomata.scala 81:44]
  wire  cam_abusy_0 = cam_s_0_state == 2'h3 | cam_amo_0; // @[AtomicAutomata.scala 82:57]
  wire  cam_dmatch_0 = cam_s_0_state != 2'h0; // @[AtomicAutomata.scala 83:49]
  wire [32:0] _a_canLogical_T_36 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_canLogical_T_38 = $signed(_a_canLogical_T_36) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  _a_canLogical_T_39 = $signed(_a_canLogical_T_38) == 33'sh0; // @[Parameters.scala 137:67]
  wire  a_isLogical = auto_in_a_bits_opcode == 3'h3; // @[AtomicAutomata.scala 90:47]
  wire  a_isArithmetic = auto_in_a_bits_opcode == 3'h2; // @[AtomicAutomata.scala 91:47]
  wire  _a_isSupported_T = a_isArithmetic ? 1'h0 : 1'h1; // @[AtomicAutomata.scala 92:63]
  wire  a_isSupported = a_isLogical ? 1'h0 : _a_isSupported_T; // @[AtomicAutomata.scala 92:32]
  wire  a_cam_busy = cam_abusy_0 & cam_a_0_fifoId == _a_canLogical_T_39; // @[AtomicAutomata.scala 105:96]
  wire  indexes_hi = cam_a_0_bits_data[0]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo = cam_d_0_data[0]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_0 = {indexes_hi,indexes_lo}; // @[Cat.scala 30:58]
  wire  indexes_hi_1 = cam_a_0_bits_data[1]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_1 = cam_d_0_data[1]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_1 = {indexes_hi_1,indexes_lo_1}; // @[Cat.scala 30:58]
  wire  indexes_hi_2 = cam_a_0_bits_data[2]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_2 = cam_d_0_data[2]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_2 = {indexes_hi_2,indexes_lo_2}; // @[Cat.scala 30:58]
  wire  indexes_hi_3 = cam_a_0_bits_data[3]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_3 = cam_d_0_data[3]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_3 = {indexes_hi_3,indexes_lo_3}; // @[Cat.scala 30:58]
  wire  indexes_hi_4 = cam_a_0_bits_data[4]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_4 = cam_d_0_data[4]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_4 = {indexes_hi_4,indexes_lo_4}; // @[Cat.scala 30:58]
  wire  indexes_hi_5 = cam_a_0_bits_data[5]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_5 = cam_d_0_data[5]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_5 = {indexes_hi_5,indexes_lo_5}; // @[Cat.scala 30:58]
  wire  indexes_hi_6 = cam_a_0_bits_data[6]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_6 = cam_d_0_data[6]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_6 = {indexes_hi_6,indexes_lo_6}; // @[Cat.scala 30:58]
  wire  indexes_hi_7 = cam_a_0_bits_data[7]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_7 = cam_d_0_data[7]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_7 = {indexes_hi_7,indexes_lo_7}; // @[Cat.scala 30:58]
  wire  indexes_hi_8 = cam_a_0_bits_data[8]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_8 = cam_d_0_data[8]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_8 = {indexes_hi_8,indexes_lo_8}; // @[Cat.scala 30:58]
  wire  indexes_hi_9 = cam_a_0_bits_data[9]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_9 = cam_d_0_data[9]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_9 = {indexes_hi_9,indexes_lo_9}; // @[Cat.scala 30:58]
  wire  indexes_hi_10 = cam_a_0_bits_data[10]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_10 = cam_d_0_data[10]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_10 = {indexes_hi_10,indexes_lo_10}; // @[Cat.scala 30:58]
  wire  indexes_hi_11 = cam_a_0_bits_data[11]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_11 = cam_d_0_data[11]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_11 = {indexes_hi_11,indexes_lo_11}; // @[Cat.scala 30:58]
  wire  indexes_hi_12 = cam_a_0_bits_data[12]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_12 = cam_d_0_data[12]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_12 = {indexes_hi_12,indexes_lo_12}; // @[Cat.scala 30:58]
  wire  indexes_hi_13 = cam_a_0_bits_data[13]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_13 = cam_d_0_data[13]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_13 = {indexes_hi_13,indexes_lo_13}; // @[Cat.scala 30:58]
  wire  indexes_hi_14 = cam_a_0_bits_data[14]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_14 = cam_d_0_data[14]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_14 = {indexes_hi_14,indexes_lo_14}; // @[Cat.scala 30:58]
  wire  indexes_hi_15 = cam_a_0_bits_data[15]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_15 = cam_d_0_data[15]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_15 = {indexes_hi_15,indexes_lo_15}; // @[Cat.scala 30:58]
  wire  indexes_hi_16 = cam_a_0_bits_data[16]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_16 = cam_d_0_data[16]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_16 = {indexes_hi_16,indexes_lo_16}; // @[Cat.scala 30:58]
  wire  indexes_hi_17 = cam_a_0_bits_data[17]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_17 = cam_d_0_data[17]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_17 = {indexes_hi_17,indexes_lo_17}; // @[Cat.scala 30:58]
  wire  indexes_hi_18 = cam_a_0_bits_data[18]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_18 = cam_d_0_data[18]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_18 = {indexes_hi_18,indexes_lo_18}; // @[Cat.scala 30:58]
  wire  indexes_hi_19 = cam_a_0_bits_data[19]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_19 = cam_d_0_data[19]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_19 = {indexes_hi_19,indexes_lo_19}; // @[Cat.scala 30:58]
  wire  indexes_hi_20 = cam_a_0_bits_data[20]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_20 = cam_d_0_data[20]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_20 = {indexes_hi_20,indexes_lo_20}; // @[Cat.scala 30:58]
  wire  indexes_hi_21 = cam_a_0_bits_data[21]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_21 = cam_d_0_data[21]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_21 = {indexes_hi_21,indexes_lo_21}; // @[Cat.scala 30:58]
  wire  indexes_hi_22 = cam_a_0_bits_data[22]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_22 = cam_d_0_data[22]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_22 = {indexes_hi_22,indexes_lo_22}; // @[Cat.scala 30:58]
  wire  indexes_hi_23 = cam_a_0_bits_data[23]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_23 = cam_d_0_data[23]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_23 = {indexes_hi_23,indexes_lo_23}; // @[Cat.scala 30:58]
  wire  indexes_hi_24 = cam_a_0_bits_data[24]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_24 = cam_d_0_data[24]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_24 = {indexes_hi_24,indexes_lo_24}; // @[Cat.scala 30:58]
  wire  indexes_hi_25 = cam_a_0_bits_data[25]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_25 = cam_d_0_data[25]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_25 = {indexes_hi_25,indexes_lo_25}; // @[Cat.scala 30:58]
  wire  indexes_hi_26 = cam_a_0_bits_data[26]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_26 = cam_d_0_data[26]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_26 = {indexes_hi_26,indexes_lo_26}; // @[Cat.scala 30:58]
  wire  indexes_hi_27 = cam_a_0_bits_data[27]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_27 = cam_d_0_data[27]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_27 = {indexes_hi_27,indexes_lo_27}; // @[Cat.scala 30:58]
  wire  indexes_hi_28 = cam_a_0_bits_data[28]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_28 = cam_d_0_data[28]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_28 = {indexes_hi_28,indexes_lo_28}; // @[Cat.scala 30:58]
  wire  indexes_hi_29 = cam_a_0_bits_data[29]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_29 = cam_d_0_data[29]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_29 = {indexes_hi_29,indexes_lo_29}; // @[Cat.scala 30:58]
  wire  indexes_hi_30 = cam_a_0_bits_data[30]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_30 = cam_d_0_data[30]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_30 = {indexes_hi_30,indexes_lo_30}; // @[Cat.scala 30:58]
  wire  indexes_hi_31 = cam_a_0_bits_data[31]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_31 = cam_d_0_data[31]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_31 = {indexes_hi_31,indexes_lo_31}; // @[Cat.scala 30:58]
  wire  indexes_hi_32 = cam_a_0_bits_data[32]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_32 = cam_d_0_data[32]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_32 = {indexes_hi_32,indexes_lo_32}; // @[Cat.scala 30:58]
  wire  indexes_hi_33 = cam_a_0_bits_data[33]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_33 = cam_d_0_data[33]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_33 = {indexes_hi_33,indexes_lo_33}; // @[Cat.scala 30:58]
  wire  indexes_hi_34 = cam_a_0_bits_data[34]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_34 = cam_d_0_data[34]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_34 = {indexes_hi_34,indexes_lo_34}; // @[Cat.scala 30:58]
  wire  indexes_hi_35 = cam_a_0_bits_data[35]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_35 = cam_d_0_data[35]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_35 = {indexes_hi_35,indexes_lo_35}; // @[Cat.scala 30:58]
  wire  indexes_hi_36 = cam_a_0_bits_data[36]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_36 = cam_d_0_data[36]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_36 = {indexes_hi_36,indexes_lo_36}; // @[Cat.scala 30:58]
  wire  indexes_hi_37 = cam_a_0_bits_data[37]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_37 = cam_d_0_data[37]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_37 = {indexes_hi_37,indexes_lo_37}; // @[Cat.scala 30:58]
  wire  indexes_hi_38 = cam_a_0_bits_data[38]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_38 = cam_d_0_data[38]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_38 = {indexes_hi_38,indexes_lo_38}; // @[Cat.scala 30:58]
  wire  indexes_hi_39 = cam_a_0_bits_data[39]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_39 = cam_d_0_data[39]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_39 = {indexes_hi_39,indexes_lo_39}; // @[Cat.scala 30:58]
  wire  indexes_hi_40 = cam_a_0_bits_data[40]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_40 = cam_d_0_data[40]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_40 = {indexes_hi_40,indexes_lo_40}; // @[Cat.scala 30:58]
  wire  indexes_hi_41 = cam_a_0_bits_data[41]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_41 = cam_d_0_data[41]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_41 = {indexes_hi_41,indexes_lo_41}; // @[Cat.scala 30:58]
  wire  indexes_hi_42 = cam_a_0_bits_data[42]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_42 = cam_d_0_data[42]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_42 = {indexes_hi_42,indexes_lo_42}; // @[Cat.scala 30:58]
  wire  indexes_hi_43 = cam_a_0_bits_data[43]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_43 = cam_d_0_data[43]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_43 = {indexes_hi_43,indexes_lo_43}; // @[Cat.scala 30:58]
  wire  indexes_hi_44 = cam_a_0_bits_data[44]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_44 = cam_d_0_data[44]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_44 = {indexes_hi_44,indexes_lo_44}; // @[Cat.scala 30:58]
  wire  indexes_hi_45 = cam_a_0_bits_data[45]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_45 = cam_d_0_data[45]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_45 = {indexes_hi_45,indexes_lo_45}; // @[Cat.scala 30:58]
  wire  indexes_hi_46 = cam_a_0_bits_data[46]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_46 = cam_d_0_data[46]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_46 = {indexes_hi_46,indexes_lo_46}; // @[Cat.scala 30:58]
  wire  indexes_hi_47 = cam_a_0_bits_data[47]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_47 = cam_d_0_data[47]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_47 = {indexes_hi_47,indexes_lo_47}; // @[Cat.scala 30:58]
  wire  indexes_hi_48 = cam_a_0_bits_data[48]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_48 = cam_d_0_data[48]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_48 = {indexes_hi_48,indexes_lo_48}; // @[Cat.scala 30:58]
  wire  indexes_hi_49 = cam_a_0_bits_data[49]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_49 = cam_d_0_data[49]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_49 = {indexes_hi_49,indexes_lo_49}; // @[Cat.scala 30:58]
  wire  indexes_hi_50 = cam_a_0_bits_data[50]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_50 = cam_d_0_data[50]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_50 = {indexes_hi_50,indexes_lo_50}; // @[Cat.scala 30:58]
  wire  indexes_hi_51 = cam_a_0_bits_data[51]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_51 = cam_d_0_data[51]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_51 = {indexes_hi_51,indexes_lo_51}; // @[Cat.scala 30:58]
  wire  indexes_hi_52 = cam_a_0_bits_data[52]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_52 = cam_d_0_data[52]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_52 = {indexes_hi_52,indexes_lo_52}; // @[Cat.scala 30:58]
  wire  indexes_hi_53 = cam_a_0_bits_data[53]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_53 = cam_d_0_data[53]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_53 = {indexes_hi_53,indexes_lo_53}; // @[Cat.scala 30:58]
  wire  indexes_hi_54 = cam_a_0_bits_data[54]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_54 = cam_d_0_data[54]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_54 = {indexes_hi_54,indexes_lo_54}; // @[Cat.scala 30:58]
  wire  indexes_hi_55 = cam_a_0_bits_data[55]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_55 = cam_d_0_data[55]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_55 = {indexes_hi_55,indexes_lo_55}; // @[Cat.scala 30:58]
  wire  indexes_hi_56 = cam_a_0_bits_data[56]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_56 = cam_d_0_data[56]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_56 = {indexes_hi_56,indexes_lo_56}; // @[Cat.scala 30:58]
  wire  indexes_hi_57 = cam_a_0_bits_data[57]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_57 = cam_d_0_data[57]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_57 = {indexes_hi_57,indexes_lo_57}; // @[Cat.scala 30:58]
  wire  indexes_hi_58 = cam_a_0_bits_data[58]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_58 = cam_d_0_data[58]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_58 = {indexes_hi_58,indexes_lo_58}; // @[Cat.scala 30:58]
  wire  indexes_hi_59 = cam_a_0_bits_data[59]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_59 = cam_d_0_data[59]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_59 = {indexes_hi_59,indexes_lo_59}; // @[Cat.scala 30:58]
  wire  indexes_hi_60 = cam_a_0_bits_data[60]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_60 = cam_d_0_data[60]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_60 = {indexes_hi_60,indexes_lo_60}; // @[Cat.scala 30:58]
  wire  indexes_hi_61 = cam_a_0_bits_data[61]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_61 = cam_d_0_data[61]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_61 = {indexes_hi_61,indexes_lo_61}; // @[Cat.scala 30:58]
  wire  indexes_hi_62 = cam_a_0_bits_data[62]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_62 = cam_d_0_data[62]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_62 = {indexes_hi_62,indexes_lo_62}; // @[Cat.scala 30:58]
  wire  indexes_hi_63 = cam_a_0_bits_data[63]; // @[AtomicAutomata.scala 113:63]
  wire  indexes_lo_63 = cam_d_0_data[63]; // @[AtomicAutomata.scala 113:73]
  wire [1:0] indexes_63 = {indexes_hi_63,indexes_lo_63}; // @[Cat.scala 30:58]
  wire [3:0] _logic_out_T = cam_a_0_lut >> indexes_0; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_lo_lo_lo_lo = _logic_out_T[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_1 = cam_a_0_lut >> indexes_1; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_lo_lo_lo_hi = _logic_out_T_1[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_2 = cam_a_0_lut >> indexes_2; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_lo_lo_hi_lo = _logic_out_T_2[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_3 = cam_a_0_lut >> indexes_3; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_lo_lo_hi_hi = _logic_out_T_3[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_4 = cam_a_0_lut >> indexes_4; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_lo_hi_lo_lo = _logic_out_T_4[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_5 = cam_a_0_lut >> indexes_5; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_lo_hi_lo_hi = _logic_out_T_5[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_6 = cam_a_0_lut >> indexes_6; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_lo_hi_hi_lo = _logic_out_T_6[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_7 = cam_a_0_lut >> indexes_7; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_lo_hi_hi_hi = _logic_out_T_7[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_8 = cam_a_0_lut >> indexes_8; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_hi_lo_lo_lo = _logic_out_T_8[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_9 = cam_a_0_lut >> indexes_9; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_hi_lo_lo_hi = _logic_out_T_9[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_10 = cam_a_0_lut >> indexes_10; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_hi_lo_hi_lo = _logic_out_T_10[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_11 = cam_a_0_lut >> indexes_11; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_hi_lo_hi_hi = _logic_out_T_11[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_12 = cam_a_0_lut >> indexes_12; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_hi_hi_lo_lo = _logic_out_T_12[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_13 = cam_a_0_lut >> indexes_13; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_hi_hi_lo_hi = _logic_out_T_13[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_14 = cam_a_0_lut >> indexes_14; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_hi_hi_hi_lo = _logic_out_T_14[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_15 = cam_a_0_lut >> indexes_15; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_lo_hi_hi_hi_hi = _logic_out_T_15[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_16 = cam_a_0_lut >> indexes_16; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_lo_lo_lo_lo = _logic_out_T_16[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_17 = cam_a_0_lut >> indexes_17; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_lo_lo_lo_hi = _logic_out_T_17[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_18 = cam_a_0_lut >> indexes_18; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_lo_lo_hi_lo = _logic_out_T_18[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_19 = cam_a_0_lut >> indexes_19; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_lo_lo_hi_hi = _logic_out_T_19[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_20 = cam_a_0_lut >> indexes_20; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_lo_hi_lo_lo = _logic_out_T_20[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_21 = cam_a_0_lut >> indexes_21; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_lo_hi_lo_hi = _logic_out_T_21[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_22 = cam_a_0_lut >> indexes_22; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_lo_hi_hi_lo = _logic_out_T_22[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_23 = cam_a_0_lut >> indexes_23; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_lo_hi_hi_hi = _logic_out_T_23[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_24 = cam_a_0_lut >> indexes_24; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_hi_lo_lo_lo = _logic_out_T_24[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_25 = cam_a_0_lut >> indexes_25; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_hi_lo_lo_hi = _logic_out_T_25[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_26 = cam_a_0_lut >> indexes_26; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_hi_lo_hi_lo = _logic_out_T_26[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_27 = cam_a_0_lut >> indexes_27; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_hi_lo_hi_hi = _logic_out_T_27[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_28 = cam_a_0_lut >> indexes_28; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_hi_hi_lo_lo = _logic_out_T_28[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_29 = cam_a_0_lut >> indexes_29; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_hi_hi_lo_hi = _logic_out_T_29[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_30 = cam_a_0_lut >> indexes_30; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_hi_hi_hi_lo = _logic_out_T_30[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_31 = cam_a_0_lut >> indexes_31; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_lo_hi_hi_hi_hi_hi = _logic_out_T_31[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_32 = cam_a_0_lut >> indexes_32; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_lo_lo_lo_lo = _logic_out_T_32[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_33 = cam_a_0_lut >> indexes_33; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_lo_lo_lo_hi = _logic_out_T_33[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_34 = cam_a_0_lut >> indexes_34; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_lo_lo_hi_lo = _logic_out_T_34[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_35 = cam_a_0_lut >> indexes_35; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_lo_lo_hi_hi = _logic_out_T_35[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_36 = cam_a_0_lut >> indexes_36; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_lo_hi_lo_lo = _logic_out_T_36[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_37 = cam_a_0_lut >> indexes_37; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_lo_hi_lo_hi = _logic_out_T_37[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_38 = cam_a_0_lut >> indexes_38; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_lo_hi_hi_lo = _logic_out_T_38[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_39 = cam_a_0_lut >> indexes_39; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_lo_hi_hi_hi = _logic_out_T_39[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_40 = cam_a_0_lut >> indexes_40; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_hi_lo_lo_lo = _logic_out_T_40[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_41 = cam_a_0_lut >> indexes_41; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_hi_lo_lo_hi = _logic_out_T_41[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_42 = cam_a_0_lut >> indexes_42; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_hi_lo_hi_lo = _logic_out_T_42[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_43 = cam_a_0_lut >> indexes_43; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_hi_lo_hi_hi = _logic_out_T_43[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_44 = cam_a_0_lut >> indexes_44; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_hi_hi_lo_lo = _logic_out_T_44[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_45 = cam_a_0_lut >> indexes_45; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_hi_hi_lo_hi = _logic_out_T_45[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_46 = cam_a_0_lut >> indexes_46; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_hi_hi_hi_lo = _logic_out_T_46[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_47 = cam_a_0_lut >> indexes_47; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_lo_hi_hi_hi_hi = _logic_out_T_47[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_48 = cam_a_0_lut >> indexes_48; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_lo_lo_lo_lo = _logic_out_T_48[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_49 = cam_a_0_lut >> indexes_49; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_lo_lo_lo_hi = _logic_out_T_49[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_50 = cam_a_0_lut >> indexes_50; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_lo_lo_hi_lo = _logic_out_T_50[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_51 = cam_a_0_lut >> indexes_51; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_lo_lo_hi_hi = _logic_out_T_51[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_52 = cam_a_0_lut >> indexes_52; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_lo_hi_lo_lo = _logic_out_T_52[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_53 = cam_a_0_lut >> indexes_53; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_lo_hi_lo_hi = _logic_out_T_53[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_54 = cam_a_0_lut >> indexes_54; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_lo_hi_hi_lo = _logic_out_T_54[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_55 = cam_a_0_lut >> indexes_55; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_lo_hi_hi_hi = _logic_out_T_55[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_56 = cam_a_0_lut >> indexes_56; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_hi_lo_lo_lo = _logic_out_T_56[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_57 = cam_a_0_lut >> indexes_57; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_hi_lo_lo_hi = _logic_out_T_57[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_58 = cam_a_0_lut >> indexes_58; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_hi_lo_hi_lo = _logic_out_T_58[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_59 = cam_a_0_lut >> indexes_59; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_hi_lo_hi_hi = _logic_out_T_59[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_60 = cam_a_0_lut >> indexes_60; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_hi_hi_lo_lo = _logic_out_T_60[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_61 = cam_a_0_lut >> indexes_61; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_hi_hi_lo_hi = _logic_out_T_61[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_62 = cam_a_0_lut >> indexes_62; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_hi_hi_hi_lo = _logic_out_T_62[0]; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_63 = cam_a_0_lut >> indexes_63; // @[AtomicAutomata.scala 114:57]
  wire  logic_out_hi_hi_hi_hi_hi_hi = _logic_out_T_63[0]; // @[AtomicAutomata.scala 114:57]
  wire [7:0] logic_out_lo_lo_lo = {logic_out_lo_lo_lo_hi_hi_hi,logic_out_lo_lo_lo_hi_hi_lo,logic_out_lo_lo_lo_hi_lo_hi,
    logic_out_lo_lo_lo_hi_lo_lo,logic_out_lo_lo_lo_lo_hi_hi,logic_out_lo_lo_lo_lo_hi_lo,logic_out_lo_lo_lo_lo_lo_hi,
    logic_out_lo_lo_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [15:0] logic_out_lo_lo = {logic_out_lo_lo_hi_hi_hi_hi,logic_out_lo_lo_hi_hi_hi_lo,logic_out_lo_lo_hi_hi_lo_hi,
    logic_out_lo_lo_hi_hi_lo_lo,logic_out_lo_lo_hi_lo_hi_hi,logic_out_lo_lo_hi_lo_hi_lo,logic_out_lo_lo_hi_lo_lo_hi,
    logic_out_lo_lo_hi_lo_lo_lo,logic_out_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] logic_out_lo_hi_lo = {logic_out_lo_hi_lo_hi_hi_hi,logic_out_lo_hi_lo_hi_hi_lo,logic_out_lo_hi_lo_hi_lo_hi,
    logic_out_lo_hi_lo_hi_lo_lo,logic_out_lo_hi_lo_lo_hi_hi,logic_out_lo_hi_lo_lo_hi_lo,logic_out_lo_hi_lo_lo_lo_hi,
    logic_out_lo_hi_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [31:0] logic_out_lo = {logic_out_lo_hi_hi_hi_hi_hi,logic_out_lo_hi_hi_hi_hi_lo,logic_out_lo_hi_hi_hi_lo_hi,
    logic_out_lo_hi_hi_hi_lo_lo,logic_out_lo_hi_hi_lo_hi_hi,logic_out_lo_hi_hi_lo_hi_lo,logic_out_lo_hi_hi_lo_lo_hi,
    logic_out_lo_hi_hi_lo_lo_lo,logic_out_lo_hi_lo,logic_out_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] logic_out_hi_lo_lo = {logic_out_hi_lo_lo_hi_hi_hi,logic_out_hi_lo_lo_hi_hi_lo,logic_out_hi_lo_lo_hi_lo_hi,
    logic_out_hi_lo_lo_hi_lo_lo,logic_out_hi_lo_lo_lo_hi_hi,logic_out_hi_lo_lo_lo_hi_lo,logic_out_hi_lo_lo_lo_lo_hi,
    logic_out_hi_lo_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [15:0] logic_out_hi_lo = {logic_out_hi_lo_hi_hi_hi_hi,logic_out_hi_lo_hi_hi_hi_lo,logic_out_hi_lo_hi_hi_lo_hi,
    logic_out_hi_lo_hi_hi_lo_lo,logic_out_hi_lo_hi_lo_hi_hi,logic_out_hi_lo_hi_lo_hi_lo,logic_out_hi_lo_hi_lo_lo_hi,
    logic_out_hi_lo_hi_lo_lo_lo,logic_out_hi_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] logic_out_hi_hi_lo = {logic_out_hi_hi_lo_hi_hi_hi,logic_out_hi_hi_lo_hi_hi_lo,logic_out_hi_hi_lo_hi_lo_hi,
    logic_out_hi_hi_lo_hi_lo_lo,logic_out_hi_hi_lo_lo_hi_hi,logic_out_hi_hi_lo_lo_hi_lo,logic_out_hi_hi_lo_lo_lo_hi,
    logic_out_hi_hi_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [31:0] logic_out_hi = {logic_out_hi_hi_hi_hi_hi_hi,logic_out_hi_hi_hi_hi_hi_lo,logic_out_hi_hi_hi_hi_lo_hi,
    logic_out_hi_hi_hi_hi_lo_lo,logic_out_hi_hi_hi_lo_hi_hi,logic_out_hi_hi_hi_lo_hi_lo,logic_out_hi_hi_hi_lo_lo_hi,
    logic_out_hi_hi_hi_lo_lo_lo,logic_out_hi_hi_lo,logic_out_hi_lo}; // @[Cat.scala 30:58]
  wire [63:0] logic_out = {logic_out_hi,logic_out_lo}; // @[Cat.scala 30:58]
  wire  unsigned_ = cam_a_0_bits_param[1]; // @[AtomicAutomata.scala 117:42]
  wire  take_max = cam_a_0_bits_param[0]; // @[AtomicAutomata.scala 118:42]
  wire  adder = cam_a_0_bits_param[2]; // @[AtomicAutomata.scala 119:39]
  wire [7:0] _signSel_T = ~cam_a_0_bits_mask; // @[AtomicAutomata.scala 121:25]
  wire [7:0] _GEN_39 = {{1'd0}, cam_a_0_bits_mask[7:1]}; // @[AtomicAutomata.scala 121:31]
  wire [7:0] _signSel_T_2 = _signSel_T | _GEN_39; // @[AtomicAutomata.scala 121:31]
  wire [7:0] signSel = ~_signSel_T_2; // @[AtomicAutomata.scala 121:23]
  wire [7:0] signbits_a = {indexes_hi_63,indexes_hi_55,indexes_hi_47,indexes_hi_39,indexes_hi_31,indexes_hi_23,
    indexes_hi_15,indexes_hi_7}; // @[Cat.scala 30:58]
  wire [7:0] signbits_d = {indexes_lo_63,indexes_lo_55,indexes_lo_47,indexes_lo_39,indexes_lo_31,indexes_lo_23,
    indexes_lo_15,indexes_lo_7}; // @[Cat.scala 30:58]
  wire [7:0] _signbit_a_T = signbits_a & signSel; // @[AtomicAutomata.scala 125:38]
  wire [8:0] _signbit_a_T_1 = {_signbit_a_T, 1'h0}; // @[AtomicAutomata.scala 125:49]
  wire [7:0] signbit_a = _signbit_a_T_1[7:0]; // @[AtomicAutomata.scala 125:54]
  wire [7:0] _signbit_d_T = signbits_d & signSel; // @[AtomicAutomata.scala 126:38]
  wire [8:0] _signbit_d_T_1 = {_signbit_d_T, 1'h0}; // @[AtomicAutomata.scala 126:49]
  wire [7:0] signbit_d = _signbit_d_T_1[7:0]; // @[AtomicAutomata.scala 126:54]
  wire [8:0] _signext_a_T = {signbit_a, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_2 = signbit_a | _signext_a_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _signext_a_T_3 = {_signext_a_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_5 = _signext_a_T_2 | _signext_a_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _signext_a_T_6 = {_signext_a_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_8 = _signext_a_T_5 | _signext_a_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] signext_a_lo_lo_lo = _signext_a_T_8[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_a_lo_lo_hi = _signext_a_T_8[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_a_lo_hi_lo = _signext_a_T_8[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_a_lo_hi_hi = _signext_a_T_8[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_a_hi_lo_lo = _signext_a_T_8[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_a_hi_lo_hi = _signext_a_T_8[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_a_hi_hi_lo = _signext_a_T_8[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_a_hi_hi_hi = _signext_a_T_8[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] signext_a = {signext_a_hi_hi_hi,signext_a_hi_hi_lo,signext_a_hi_lo_hi,signext_a_hi_lo_lo,
    signext_a_lo_hi_hi,signext_a_lo_hi_lo,signext_a_lo_lo_hi,signext_a_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [8:0] _signext_d_T = {signbit_d, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_2 = signbit_d | _signext_d_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _signext_d_T_3 = {_signext_d_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_5 = _signext_d_T_2 | _signext_d_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _signext_d_T_6 = {_signext_d_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_8 = _signext_d_T_5 | _signext_d_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] signext_d_lo_lo_lo = _signext_d_T_8[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_d_lo_lo_hi = _signext_d_T_8[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_d_lo_hi_lo = _signext_d_T_8[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_d_lo_hi_hi = _signext_d_T_8[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_d_hi_lo_lo = _signext_d_T_8[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_d_hi_lo_hi = _signext_d_T_8[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_d_hi_hi_lo = _signext_d_T_8[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] signext_d_hi_hi_hi = _signext_d_T_8[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] signext_d = {signext_d_hi_hi_hi,signext_d_hi_hi_lo,signext_d_hi_lo_hi,signext_d_hi_lo_lo,
    signext_d_lo_hi_hi,signext_d_lo_hi_lo,signext_d_lo_lo_hi,signext_d_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] wide_mask_lo_lo_lo = cam_a_0_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] wide_mask_lo_lo_hi = cam_a_0_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] wide_mask_lo_hi_lo = cam_a_0_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] wide_mask_lo_hi_hi = cam_a_0_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] wide_mask_hi_lo_lo = cam_a_0_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] wide_mask_hi_lo_hi = cam_a_0_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] wide_mask_hi_hi_lo = cam_a_0_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] wide_mask_hi_hi_hi = cam_a_0_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] wide_mask = {wide_mask_hi_hi_hi,wide_mask_hi_hi_lo,wide_mask_hi_lo_hi,wide_mask_hi_lo_lo,
    wide_mask_lo_hi_hi,wide_mask_lo_hi_lo,wide_mask_lo_lo_hi,wide_mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _a_a_ext_T = cam_a_0_bits_data & wide_mask; // @[AtomicAutomata.scala 131:28]
  wire [63:0] a_a_ext = _a_a_ext_T | signext_a; // @[AtomicAutomata.scala 131:41]
  wire [63:0] _a_d_ext_T = cam_d_0_data & wide_mask; // @[AtomicAutomata.scala 132:28]
  wire [63:0] a_d_ext = _a_d_ext_T | signext_d; // @[AtomicAutomata.scala 132:41]
  wire [63:0] _a_d_inv_T = ~a_d_ext; // @[AtomicAutomata.scala 133:43]
  wire [63:0] a_d_inv = adder ? a_d_ext : _a_d_inv_T; // @[AtomicAutomata.scala 133:26]
  wire [63:0] adder_out = a_a_ext + a_d_inv; // @[AtomicAutomata.scala 134:33]
  wire  a_bigger_uneq = unsigned_ == a_a_ext[63]; // @[AtomicAutomata.scala 136:38]
  wire  a_bigger = a_a_ext[63] == a_d_ext[63] ? ~adder_out[63] : a_bigger_uneq; // @[AtomicAutomata.scala 137:27]
  wire  pick_a = take_max == a_bigger; // @[AtomicAutomata.scala 138:31]
  wire [63:0] _arith_out_T = pick_a ? cam_a_0_bits_data : cam_d_0_data; // @[AtomicAutomata.scala 139:50]
  wire [63:0] arith_out = adder ? adder_out : _arith_out_T; // @[AtomicAutomata.scala 139:28]
  wire [63:0] amo_data = cam_a_0_bits_opcode[0] ? logic_out : arith_out; // @[AtomicAutomata.scala 145:14]
  wire  a_allow = ~a_cam_busy & (a_isSupported | cam_free_0); // @[AtomicAutomata.scala 149:35]
  reg [2:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 3'h0; // @[Arbiter.scala 88:28]
  wire  source_i_valid = auto_in_a_valid & a_allow; // @[AtomicAutomata.scala 151:38]
  wire [1:0] _readys_T = {source_i_valid,cam_amo_0}; // @[Cat.scala 30:58]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[package.scala 244:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[Arbiter.scala 16:61]
  wire  readys_1 = _readys_T_7[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 123:31]
  wire  _T = ~a_isSupported; // @[AtomicAutomata.scala 153:15]
  wire [2:0] source_i_bits_opcode = ~a_isSupported ? 3'h4 : auto_in_a_bits_opcode; // @[AtomicAutomata.scala 153:31 AtomicAutomata.scala 154:32 AtomicAutomata.scala 152:24]
  wire [2:0] source_i_bits_param = ~a_isSupported ? 3'h0 : auto_in_a_bits_param; // @[AtomicAutomata.scala 153:31 AtomicAutomata.scala 155:32 AtomicAutomata.scala 152:24]
  wire [1:0] source_c_bits_a_mask_sizeOH_shiftAmount = cam_a_0_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _source_c_bits_a_mask_sizeOH_T_1 = 4'h1 << source_c_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] source_c_bits_a_mask_sizeOH = _source_c_bits_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _source_c_bits_a_mask_T = cam_a_0_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  source_c_bits_a_mask_size = source_c_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit = cam_a_0_bits_address[2]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit = ~source_c_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_acc = _source_c_bits_a_mask_T | source_c_bits_a_mask_size & source_c_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_acc_1 = _source_c_bits_a_mask_T | source_c_bits_a_mask_size & source_c_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_size_1 = source_c_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit_1 = cam_a_0_bits_address[1]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit_1 = ~source_c_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_eq_2 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_2 = source_c_bits_a_mask_acc | source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_3 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_3 = source_c_bits_a_mask_acc | source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_4 = source_c_bits_a_mask_bit & source_c_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_4 = source_c_bits_a_mask_acc_1 | source_c_bits_a_mask_size_1 &
    source_c_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_5 = source_c_bits_a_mask_bit & source_c_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_5 = source_c_bits_a_mask_acc_1 | source_c_bits_a_mask_size_1 &
    source_c_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_size_2 = source_c_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit_2 = cam_a_0_bits_address[0]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit_2 = ~source_c_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_eq_6 = source_c_bits_a_mask_eq_2 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_lo_lo_lo = source_c_bits_a_mask_acc_2 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_7 = source_c_bits_a_mask_eq_2 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_lo_lo_hi = source_c_bits_a_mask_acc_2 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_8 = source_c_bits_a_mask_eq_3 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_lo_hi_lo = source_c_bits_a_mask_acc_3 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_9 = source_c_bits_a_mask_eq_3 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_lo_hi_hi = source_c_bits_a_mask_acc_3 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_10 = source_c_bits_a_mask_eq_4 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_hi_lo_lo = source_c_bits_a_mask_acc_4 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_11 = source_c_bits_a_mask_eq_4 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_hi_lo_hi = source_c_bits_a_mask_acc_4 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_12 = source_c_bits_a_mask_eq_5 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_hi_hi_lo = source_c_bits_a_mask_acc_5 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_13 = source_c_bits_a_mask_eq_5 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_hi_hi_hi = source_c_bits_a_mask_acc_5 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] source_c_bits_a_mask = {source_c_bits_a_mask_hi_hi_hi,source_c_bits_a_mask_hi_hi_lo,
    source_c_bits_a_mask_hi_lo_hi,source_c_bits_a_mask_hi_lo_lo,source_c_bits_a_mask_lo_hi_hi,
    source_c_bits_a_mask_lo_hi_lo,source_c_bits_a_mask_lo_lo_hi,source_c_bits_a_mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [12:0] _decode_T_1 = 13'h3f << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _decode_T_3 = ~_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] decode = _decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 89:24]
  wire  readys_0 = _readys_T_7[0]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_0 = readys_0 & cam_amo_0; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1 = readys_1 & source_i_valid; // @[Arbiter.scala 97:79]
  wire  _prefixOR_T = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 104:53]
  wire  _T_12 = cam_amo_0 | source_i_valid; // @[Arbiter.scala 107:36]
  wire  _T_13 = ~(cam_amo_0 | source_i_valid); // @[Arbiter.scala 107:15]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & cam_amo_0 | state_1 & source_i_valid; // @[Mux.scala 27:72]
  wire  sink_ACancel_earlyValid = idle ? _T_12 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 50:33]
  wire [2:0] _GEN_40 = {{2'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [2:0] _beatsLeft_T_4 = beatsLeft - _GEN_40; // @[Arbiter.scala 113:52]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  out_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  wire [63:0] _T_29 = muxStateEarly_0 ? amo_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_30 = muxStateEarly_1 ? auto_in_a_bits_data : 64'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_32 = muxStateEarly_0 ? source_c_bits_a_mask : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_33 = muxStateEarly_1 ? auto_in_a_bits_mask : 8'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_35 = muxStateEarly_0 ? cam_a_0_bits_address : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_36 = muxStateEarly_1 ? auto_in_a_bits_address : 32'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_38 = muxStateEarly_0 ? cam_a_0_bits_source : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_39 = muxStateEarly_1 ? auto_in_a_bits_source : 7'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_41 = muxStateEarly_0 ? cam_a_0_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_42 = muxStateEarly_1 ? auto_in_a_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire  _T_50 = out_1_ready & source_i_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_41 = {{1'd0}, auto_in_a_bits_param[1:0]}; // @[Mux.scala 80:60]
  wire [3:0] _cam_a_0_lut_T_2 = 3'h1 == _GEN_41 ? 4'he : 4'h8; // @[Mux.scala 80:57]
  wire [1:0] _GEN_12 = cam_free_0 ? 2'h3 : cam_s_0_state; // @[AtomicAutomata.scala 187:23 AtomicAutomata.scala 188:23 AtomicAutomata.scala 76:28]
  wire [1:0] _GEN_23 = _T_50 & _T ? _GEN_12 : cam_s_0_state; // @[AtomicAutomata.scala 174:50 AtomicAutomata.scala 76:28]
  wire  _T_53 = out_ready & cam_amo_0; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_24 = cam_amo_0 ? 2'h1 : _GEN_23; // @[AtomicAutomata.scala 196:23 AtomicAutomata.scala 197:23]
  wire [1:0] _GEN_25 = _T_53 ? _GEN_24 : _GEN_23; // @[AtomicAutomata.scala 194:32]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  wire  d_ackd = auto_out_d_bits_opcode == 3'h1; // @[AtomicAutomata.scala 213:40]
  wire  d_cam_sel_raw_0 = cam_a_0_bits_source == auto_out_d_bits_source; // @[AtomicAutomata.scala 204:53]
  wire  d_cam_sel_match_0 = d_cam_sel_raw_0 & cam_dmatch_0; // @[AtomicAutomata.scala 205:83]
  wire  d_drop = d_first & d_ackd & d_cam_sel_match_0; // @[AtomicAutomata.scala 232:40]
  wire  bundleOut_0_d_ready = auto_in_d_ready | d_drop; // @[AtomicAutomata.scala 236:35]
  wire  _d_first_T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_ack = auto_out_d_bits_opcode == 3'h0; // @[AtomicAutomata.scala 214:40]
  wire  d_replace = d_first & d_ack & d_cam_sel_match_0; // @[AtomicAutomata.scala 233:42]
  TLMonitor_12 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_c_ready(monitor_io_in_c_ready),
    .io_in_c_valid(monitor_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_io_in_c_bits_address),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),
    .io_in_e_ready(monitor_io_in_e_ready),
    .io_in_e_valid(monitor_io_in_e_valid),
    .io_in_e_bits_sink(monitor_io_in_e_bits_sink)
  );
  assign auto_in_a_ready = out_1_ready & a_allow; // @[AtomicAutomata.scala 150:38]
  assign auto_in_c_ready = auto_out_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_valid = auto_out_d_valid & ~d_drop; // @[AtomicAutomata.scala 235:35]
  assign auto_in_d_bits_opcode = d_replace ? 3'h1 : auto_out_d_bits_opcode; // @[AtomicAutomata.scala 239:26 AtomicAutomata.scala 240:28 AtomicAutomata.scala 238:19]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = d_replace ? cam_d_0_denied | auto_out_d_bits_denied : auto_out_d_bits_denied; // @[AtomicAutomata.scala 239:26 AtomicAutomata.scala 243:29 AtomicAutomata.scala 238:19]
  assign auto_in_d_bits_data = d_replace ? cam_d_0_data : auto_out_d_bits_data; // @[AtomicAutomata.scala 239:26 AtomicAutomata.scala 241:26 AtomicAutomata.scala 238:19]
  assign auto_in_d_bits_corrupt = d_replace ? cam_d_0_corrupt | auto_out_d_bits_denied : auto_out_d_bits_corrupt; // @[AtomicAutomata.scala 239:26 AtomicAutomata.scala 242:29 AtomicAutomata.scala 238:19]
  assign auto_in_e_ready = auto_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = idle ? _T_12 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_out_a_bits_opcode = muxStateEarly_1 ? source_i_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  assign auto_out_a_bits_param = muxStateEarly_1 ? source_i_bits_param : 3'h0; // @[Mux.scala 27:72]
  assign auto_out_a_bits_size = _T_41 | _T_42; // @[Mux.scala 27:72]
  assign auto_out_a_bits_source = _T_38 | _T_39; // @[Mux.scala 27:72]
  assign auto_out_a_bits_address = _T_35 | _T_36; // @[Mux.scala 27:72]
  assign auto_out_a_bits_mask = _T_32 | _T_33; // @[Mux.scala 27:72]
  assign auto_out_a_bits_data = _T_29 | _T_30; // @[Mux.scala 27:72]
  assign auto_out_a_bits_corrupt = muxStateEarly_0 & cam_d_0_corrupt; // @[Mux.scala 27:72]
  assign auto_out_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready | d_drop; // @[AtomicAutomata.scala 236:35]
  assign auto_out_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = out_1_ready & a_allow; // @[AtomicAutomata.scala 150:38]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_ready = auto_out_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = auto_out_d_valid & ~d_drop; // @[AtomicAutomata.scala 235:35]
  assign monitor_io_in_d_bits_opcode = d_replace ? 3'h1 : auto_out_d_bits_opcode; // @[AtomicAutomata.scala 239:26 AtomicAutomata.scala 240:28 AtomicAutomata.scala 238:19]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_denied = d_replace ? cam_d_0_denied | auto_out_d_bits_denied : auto_out_d_bits_denied; // @[AtomicAutomata.scala 239:26 AtomicAutomata.scala 243:29 AtomicAutomata.scala 238:19]
  assign monitor_io_in_d_bits_corrupt = d_replace ? cam_d_0_corrupt | auto_out_d_bits_denied : auto_out_d_bits_corrupt; // @[AtomicAutomata.scala 239:26 AtomicAutomata.scala 242:29 AtomicAutomata.scala 238:19]
  assign monitor_io_in_e_ready = auto_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  always @(posedge clock) begin
    if (reset) begin // @[AtomicAutomata.scala 76:28]
      cam_s_0_state <= 2'h0; // @[AtomicAutomata.scala 76:28]
    end else if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0) begin // @[AtomicAutomata.scala 225:23]
        if (d_ackd) begin // @[AtomicAutomata.scala 227:29]
          cam_s_0_state <= 2'h2;
        end else begin
          cam_s_0_state <= 2'h0;
        end
      end else begin
        cam_s_0_state <= _GEN_25;
      end
    end else begin
      cam_s_0_state <= _GEN_25;
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        cam_a_0_bits_opcode <= auto_in_a_bits_opcode; // @[AtomicAutomata.scala 178:24]
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        cam_a_0_bits_param <= auto_in_a_bits_param; // @[AtomicAutomata.scala 178:24]
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        cam_a_0_bits_size <= auto_in_a_bits_size; // @[AtomicAutomata.scala 178:24]
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        cam_a_0_bits_source <= auto_in_a_bits_source; // @[AtomicAutomata.scala 178:24]
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        cam_a_0_bits_address <= auto_in_a_bits_address; // @[AtomicAutomata.scala 178:24]
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        cam_a_0_bits_mask <= auto_in_a_bits_mask; // @[AtomicAutomata.scala 178:24]
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        cam_a_0_bits_data <= auto_in_a_bits_data; // @[AtomicAutomata.scala 178:24]
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        cam_a_0_fifoId <= _a_canLogical_T_39; // @[AtomicAutomata.scala 177:24]
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin // @[AtomicAutomata.scala 176:23]
        if (3'h3 == _GEN_41) begin // @[Mux.scala 80:57]
          cam_a_0_lut <= 4'hc;
        end else if (3'h0 == _GEN_41) begin // @[Mux.scala 80:57]
          cam_a_0_lut <= 4'h6;
        end else begin
          cam_a_0_lut <= _cam_a_0_lut_T_2;
        end
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin // @[AtomicAutomata.scala 218:33]
        cam_d_0_data <= auto_out_d_bits_data; // @[AtomicAutomata.scala 219:22]
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin // @[AtomicAutomata.scala 218:33]
        cam_d_0_denied <= auto_out_d_bits_denied; // @[AtomicAutomata.scala 220:24]
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin // @[AtomicAutomata.scala 218:33]
        cam_d_0_corrupt <= auto_out_d_bits_corrupt; // @[AtomicAutomata.scala 221:25]
      end
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 3'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin // @[Arbiter.scala 113:23]
      if (earlyWinner_1) begin // @[Arbiter.scala 111:73]
        if (opdata) begin // @[Edges.scala 220:14]
          beatsLeft <= decode;
        end else begin
          beatsLeft <= 3'h0;
        end
      end else begin
        beatsLeft <= 3'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin // @[Arbiter.scala 117:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin // @[Arbiter.scala 117:30]
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1 | reset)) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(cam_amo_0 | source_i_valid) | _prefixOR_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(cam_amo_0 | source_i_valid) | _prefixOR_T | reset)) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_13 | _T_12 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_13 | _T_12 | reset)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cam_s_0_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cam_a_0_bits_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  cam_a_0_bits_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  cam_a_0_bits_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  cam_a_0_bits_source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  cam_a_0_bits_address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cam_a_0_bits_mask = _RAND_6[7:0];
  _RAND_7 = {2{`RANDOM}};
  cam_a_0_bits_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  cam_a_0_fifoId = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  cam_a_0_lut = _RAND_9[3:0];
  _RAND_10 = {2{`RANDOM}};
  cam_d_0_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  cam_d_0_denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  cam_d_0_corrupt = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  beatsLeft = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  state_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  d_first_counter = _RAND_16[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_13(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [2:0]  io_in_c_bits_size,
  input  [6:0]  io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [6:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input         io_in_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_86 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_2 = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_3 = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_4 = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_5 = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_lo = mask_acc_2 | mask_size_2 & mask_eq_6; // @[Misc.scala 214:29]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_hi = mask_acc_2 | mask_size_2 & mask_eq_7; // @[Misc.scala 214:29]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_lo = mask_acc_3 | mask_size_2 & mask_eq_8; // @[Misc.scala 214:29]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_hi = mask_acc_3 | mask_size_2 & mask_eq_9; // @[Misc.scala 214:29]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_lo = mask_acc_4 | mask_size_2 & mask_eq_10; // @[Misc.scala 214:29]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_hi = mask_acc_4 | mask_size_2 & mask_eq_11; // @[Misc.scala 214:29]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_lo = mask_acc_5 | mask_size_2 & mask_eq_12; // @[Misc.scala 214:29]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_hi = mask_acc_5 | mask_size_2 & mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire [31:0] _T_180 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_181 = {1'b0,$signed(_T_180)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_183 = $signed(_T_181) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_184 = $signed(_T_183) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_185 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_186 = {1'b0,$signed(_T_185)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_188 = $signed(_T_186) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_189 = $signed(_T_188) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_190 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_191 = {1'b0,$signed(_T_190)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_193 = $signed(_T_191) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_194 = $signed(_T_193) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_195 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_196 = {1'b0,$signed(_T_195)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_198 = $signed(_T_196) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_199 = $signed(_T_198) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_200 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_201 = {1'b0,$signed(_T_200)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_203 = $signed(_T_201) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_204 = $signed(_T_203) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_211 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_214 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_215 = {1'b0,$signed(_T_214)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_217 = $signed(_T_215) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_218 = $signed(_T_217) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_219 = _T_211 & _T_218; // @[Parameters.scala 670:56]
  wire  _T_222 = source_ok & _T_219; // @[Monitor.scala 82:72]
  wire  _T_277 = _source_ok_T_1 & _T_211; // @[Mux.scala 27:72]
  wire  _T_330 = _T_218 | _T_184 | _T_189 | _T_194 | _T_199 | _T_204; // @[Parameters.scala 671:42]
  wire  _T_333 = _T_277 & _T_330; // @[Monitor.scala 83:78]
  wire  _T_347 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [7:0] _T_351 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_352 = _T_351 == 8'h0; // @[Monitor.scala 88:31]
  wire  _T_360 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_593 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_606 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_709 = _T_211 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_720 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_724 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_732 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_834 = source_ok & _T_709; // @[Monitor.scala 115:71]
  wire  _T_852 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [7:0] _T_968 = ~mask; // @[Monitor.scala 127:33]
  wire [7:0] _T_969 = io_in_a_bits_mask & _T_968; // @[Monitor.scala 127:31]
  wire  _T_970 = _T_969 == 8'h0; // @[Monitor.scala 127:40]
  wire  _T_974 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_1036 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_1074 = _T_1036 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_1076 = source_ok & _T_1074; // @[Monitor.scala 131:74]
  wire  _T_1086 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_1094 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_1206 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_1214 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1328 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1340 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1344 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1348 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27]
  wire  _T_1352 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_1356 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1360 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1364 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1375 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_1379 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_1392 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1412 = _T_1360 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1421 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1438 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1456 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _source_ok_T_109 = io_in_c_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_115 = io_in_c_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_121 = io_in_c_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_127 = io_in_c_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_133 = io_in_c_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_139 = io_in_c_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_145 = io_in_c_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_151 = io_in_c_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_2 = _source_ok_T_109 | _source_ok_T_115 | _source_ok_T_121 | _source_ok_T_127 | _source_ok_T_133 |
    _source_ok_T_139 | _source_ok_T_145 | _source_ok_T_151; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_7 = 13'h3f << io_in_c_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask_2 = ~_is_aligned_mask_T_7[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_87 = {{26'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T_2 = io_in_c_bits_address & _GEN_87; // @[Edges.scala 20:16]
  wire  is_aligned_2 = _is_aligned_T_2 == 32'h0; // @[Edges.scala 20:24]
  wire [31:0] _address_ok_T_34 = io_in_c_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_35 = {1'b0,$signed(_address_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_37 = $signed(_address_ok_T_35) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_38 = $signed(_address_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_39 = io_in_c_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_40 = {1'b0,$signed(_address_ok_T_39)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_42 = $signed(_address_ok_T_40) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_43 = $signed(_address_ok_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_44 = io_in_c_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_45 = {1'b0,$signed(_address_ok_T_44)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_47 = $signed(_address_ok_T_45) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_48 = $signed(_address_ok_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_49 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_50 = {1'b0,$signed(_address_ok_T_49)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_52 = $signed(_address_ok_T_50) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_53 = $signed(_address_ok_T_52) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_54 = io_in_c_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_55 = {1'b0,$signed(_address_ok_T_54)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_57 = $signed(_address_ok_T_55) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_58 = $signed(_address_ok_T_57) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _address_ok_T_62 = _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 | _address_ok_T_58; // @[Parameters.scala 598:92]
  wire [31:0] _address_ok_T_63 = io_in_c_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_64 = {1'b0,$signed(_address_ok_T_63)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_66 = $signed(_address_ok_T_64) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_67 = $signed(_address_ok_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  wire  address_ok_1 = _address_ok_T_62 | _address_ok_T_67; // @[Parameters.scala 622:64]
  wire  _T_2226 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  wire  _T_2233 = io_in_c_bits_size >= 3'h3; // @[Monitor.scala 245:30]
  wire  _T_2240 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  wire  _T_2248 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  wire  _T_2266 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  wire  _T_2359 = io_in_c_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_2367 = _T_2359 & _address_ok_T_67; // @[Parameters.scala 670:56]
  wire  _T_2370 = source_ok_2 & _T_2367; // @[Monitor.scala 260:78]
  wire  _T_2425 = _source_ok_T_109 & _T_2359; // @[Mux.scala 27:72]
  wire  _T_2478 = _address_ok_T_67 | _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 |
    _address_ok_T_58; // @[Parameters.scala 671:42]
  wire  _T_2481 = _T_2425 & _T_2478; // @[Monitor.scala 261:78]
  wire  _T_2503 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  wire  _T_2736 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  wire  _T_2746 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  wire  _T_2754 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  wire  _T_2768 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  wire  sink_ok_1 = io_in_e_bits_sink < 1'h1; // @[Monitor.scala 364:31]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [6:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_2790 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_2791 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_2795 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_2799 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_2803 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_2807 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [6:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_2814 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_2815 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_2819 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_2823 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_2827 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_2835 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  wire  _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  wire [2:0] c_first_beats1_decode = is_aligned_mask_2[5:3]; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  reg [2:0] c_first_counter; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1 = c_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  c_first = c_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [2:0] size_3; // @[Monitor.scala 514:22]
  reg [6:0] source_3; // @[Monitor.scala 515:22]
  reg [31:0] address_2; // @[Monitor.scala 516:22]
  wire  _T_2866 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  wire  _T_2867 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  wire  _T_2871 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  wire  _T_2875 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  wire  _T_2879 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  wire  _T_2883 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  reg [127:0] inflight; // @[Monitor.scala 611:27]
  reg [511:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [511:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  wire [8:0] _GEN_88 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [9:0] _a_opcode_lookup_T = {{1'd0}, _GEN_88}; // @[Monitor.scala 634:69]
  wire [511:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [511:0] _GEN_89 = {{496'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_89; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[511:1]}; // @[Monitor.scala 634:152]
  wire [511:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [511:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 638:91]
  wire [511:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[511:1]}; // @[Monitor.scala 638:144]
  wire  _T_2889 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [127:0] _a_set_wo_ready_T = 128'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_2892 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [8:0] _GEN_94 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [9:0] _a_opcodes_set_T = {{1'd0}, _GEN_94}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [1026:0] _GEN_95 = {{1023'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [1026:0] _a_opcodes_set_T_1 = _GEN_95 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [1026:0] _GEN_97 = {{1023'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [1026:0] _a_sizes_set_T_1 = _GEN_97 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [127:0] _T_2894 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_2896 = ~_T_2894[0]; // @[Monitor.scala 658:17]
  wire [127:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [1026:0] _GEN_31 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [1026:0] _GEN_32 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_2900 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_2902 = ~_T_1344; // @[Monitor.scala 671:74]
  wire  _T_2903 = io_in_d_valid & d_first_1 & ~_T_1344; // @[Monitor.scala 671:71]
  wire [127:0] _d_clr_wo_ready_T = 128'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1344 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [1038:0] _GEN_99 = {{1023'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [1038:0] _d_opcodes_clr_T_5 = _GEN_99 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [127:0] d_clr = _d_first_T & d_first_1 & _T_2902 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [1038:0] _GEN_35 = _d_first_T & d_first_1 & _T_2902 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_2889 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [127:0] _T_2913 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_2915 = _T_2913[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_2920 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_2921 = io_in_d_bits_opcode == _GEN_44 | _T_2920; // @[Monitor.scala 685:77]
  wire  _T_2925 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_2932 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_2933 = io_in_d_bits_opcode == _GEN_60 | _T_2932; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_102 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_2937 = _GEN_102 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_2947 = _T_2900 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_2902; // @[Monitor.scala 694:116]
  wire  _T_2948 = ~io_in_d_ready; // @[Monitor.scala 695:15]
  wire  _T_2949 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_2956 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [127:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [127:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [127:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [511:0] a_opcodes_set = _GEN_31[511:0];
  wire [511:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [511:0] d_opcodes_clr = _GEN_35[511:0];
  wire [511:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [511:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [511:0] a_sizes_set = _GEN_32[511:0];
  wire [511:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [511:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_2965 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [127:0] inflight_1; // @[Monitor.scala 723:35]
  reg [511:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [2:0] c_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1_1 = c_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  c_first_1 = c_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25]
  wire [511:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [511:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 747:93]
  wire [511:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[511:1]}; // @[Monitor.scala 747:146]
  wire  _T_2975 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  _T_2976 = io_in_c_valid & c_first_1 & _T_2975; // @[Monitor.scala 756:37]
  wire [127:0] _c_set_wo_ready_T = 128'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] c_set_wo_ready = io_in_c_valid & c_first_1 & _T_2975 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 756:71 Monitor.scala 757:22]
  wire  _T_2982 = _c_first_T & c_first_1 & _T_2975; // @[Monitor.scala 760:38]
  wire [3:0] _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  wire [3:0] _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 4'h1; // @[Monitor.scala 763:59]
  wire [8:0] _GEN_109 = {io_in_c_bits_source, 2'h0}; // @[Monitor.scala 764:79]
  wire [9:0] _c_opcodes_set_T = {{1'd0}, _GEN_109}; // @[Monitor.scala 764:79]
  wire [3:0] c_sizes_set_interm = _c_first_T & c_first_1 & _T_2975 ? _c_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 760:72 Monitor.scala 763:28]
  wire [1026:0] _GEN_112 = {{1023'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  wire [1026:0] _c_sizes_set_T_1 = _GEN_112 << _c_opcodes_set_T; // @[Monitor.scala 765:52]
  wire [127:0] _T_2983 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  wire  _T_2985 = ~_T_2983[0]; // @[Monitor.scala 766:17]
  wire [127:0] c_set = _c_first_T & c_first_1 & _T_2975 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 760:72 Monitor.scala 761:28]
  wire [1026:0] _GEN_77 = _c_first_T & c_first_1 & _T_2975 ? _c_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 760:72 Monitor.scala 765:28]
  wire  _T_2989 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  wire  _T_2991 = io_in_d_valid & d_first_2 & _T_1344; // @[Monitor.scala 779:71]
  wire [127:0] d_clr_wo_ready_1 = io_in_d_valid & d_first_2 & _T_1344 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 779:89 Monitor.scala 780:22]
  wire [127:0] d_clr_1 = _d_first_T & d_first_2 & _T_1344 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [1038:0] _GEN_80 = _d_first_T & d_first_2 & _T_1344 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire  _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1 = _T_2976 & io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:88]
  wire [127:0] _T_2999 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire  _T_3001 = _T_2999[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  wire  _T_3005 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_3009 = _GEN_102 == c_size_lookup; // @[Monitor.scala 795:36]
  wire  _T_3018 = _T_2989 & c_first_1 & io_in_c_valid & _same_cycle_resp_T_8 & _T_1344; // @[Monitor.scala 799:116]
  wire  _T_3020 = _T_2948 | io_in_c_ready; // @[Monitor.scala 800:32]
  wire  _T_3024 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  wire  _T_3025 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  wire [127:0] _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  wire [127:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [127:0] _inflight_T_5 = _inflight_T_3 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [511:0] d_opcodes_clr_1 = _GEN_80[511:0];
  wire [511:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [511:0] c_sizes_set = _GEN_77[511:0];
  wire [511:0] _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  wire [511:0] _inflight_sizes_T_5 = _inflight_sizes_T_3 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_3034 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [2:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_3 = d_first_counter_3 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 3'h0; // @[Edges.scala 230:25]
  wire  _T_3046 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_3047 = _d_first_T & d_first_3 & _T_3046; // @[Monitor.scala 829:38]
  wire  _T_3050 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = _d_first_T & d_first_3 & _T_3046 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  _T_3054 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _e_clr_T = 2'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  wire  d_set = _GEN_84[0];
  wire  _T_3058 = (d_set | inflight_2) >> io_in_e_bits_sink; // @[Monitor.scala 837:35]
  wire [1:0] _GEN_85 = _T_3054 ? _e_clr_T : 2'h0; // @[Monitor.scala 835:73 Monitor.scala 836:13]
  wire  e_clr = _GEN_85[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 3'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      opcode_3 <= io_in_c_bits_opcode; // @[Monitor.scala 525:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      param_3 <= io_in_c_bits_param; // @[Monitor.scala 526:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      size_3 <= io_in_c_bits_size; // @[Monitor.scala 527:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      source_3 <= io_in_c_bits_source; // @[Monitor.scala 528:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      address_2 <= io_in_c_bits_address; // @[Monitor.scala 529:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 128'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 512'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 512'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 128'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 512'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first_1) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 3'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_c_first_T | _d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= (inflight_2 | d_set) & ~e_clr; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 3'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1328 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1328 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1340 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1340 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1348 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1348 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1360 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1344 & ~(_T_1360 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1348 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1348 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1375 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1375 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1379 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1379 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1364 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1348 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1348 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1375 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1375 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1379 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1379 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1412 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1392 & ~(_T_1412 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1421 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(_T_1412 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1438 & ~(_T_1412 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(_T_1352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(_T_1352 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(_T_1356 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1456 & ~(_T_1356 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(_T_2233 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(_T_2233 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(_T_2240 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2226 & ~(_T_2240 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(_T_2233 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(_T_2233 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(_T_2240 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2248 & ~(_T_2240 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2370 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2370 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2481 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2481 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2233 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2233 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2240 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid report param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2266 & ~(_T_2240 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2370 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2370 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2481 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2481 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2233 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2233 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2240 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2503 & ~(_T_2240 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(_T_2746 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2736 & ~(_T_2746 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(_T_2746 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2754 & ~(_T_2746 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(_T_2746 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2768 & ~(_T_2746 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channels carries invalid sink ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2791 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2791 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2795 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2795 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2799 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2799 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2803 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2803 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2790 & ~(_T_2807 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2790 & ~(_T_2807 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2815 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2815 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2819 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2819 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2823 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2823 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2827 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2827 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2814 & ~(_T_2835 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2814 & ~(_T_2835 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2867 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2867 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2871 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2871 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2875 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2875 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2879 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2879 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2866 & ~(_T_2883 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2866 & ~(_T_2883 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2892 & ~(_T_2896 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2892 & ~(_T_2896 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & ~(_T_2915 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & ~(_T_2915 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & same_cycle_resp & ~(_T_2921 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & same_cycle_resp & ~(_T_2921 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & same_cycle_resp & ~(_T_2925 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & same_cycle_resp & ~(_T_2925 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & ~same_cycle_resp & ~(_T_2933 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & ~same_cycle_resp & ~(_T_2933 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2903 & ~same_cycle_resp & ~(_T_2937 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2903 & ~same_cycle_resp & ~(_T_2937 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2947 & ~(_T_2949 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2947 & ~(_T_2949 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2956 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2956 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2965 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2965 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2982 & ~(_T_2985 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel re-used a source ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2982 & ~(_T_2985 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2991 & ~(_T_3001 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2991 & ~(_T_3001 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2991 & same_cycle_resp_1 & ~(_T_3005 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2991 & same_cycle_resp_1 & ~(_T_3005 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2991 & ~same_cycle_resp_1 & ~(_T_3009 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2991 & ~same_cycle_resp_1 & ~(_T_3009 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3018 & ~(_T_3020 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3018 & ~(_T_3020 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3024 & ~(_T_3025 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3024 & ~(_T_3025 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_3034 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_3034 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3047 & ~(_T_3050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3047 & ~(_T_3050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3054 & ~(_T_3058 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:79)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3054 & ~(_T_3058 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  c_first_counter = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  opcode_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  param_3 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  size_3 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  source_3 = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  address_2 = _RAND_17[31:0];
  _RAND_18 = {4{`RANDOM}};
  inflight = _RAND_18[127:0];
  _RAND_19 = {16{`RANDOM}};
  inflight_opcodes = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  inflight_sizes = _RAND_20[511:0];
  _RAND_21 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  watchdog = _RAND_23[31:0];
  _RAND_24 = {4{`RANDOM}};
  inflight_1 = _RAND_24[127:0];
  _RAND_25 = {16{`RANDOM}};
  inflight_sizes_1 = _RAND_25[511:0];
  _RAND_26 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  watchdog_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inflight_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_30[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFIFOFixer_1(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [2:0]  auto_in_c_bits_size,
  input  [6:0]  auto_in_c_bits_source,
  input  [31:0] auto_in_c_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  output        auto_in_e_ready,
  input         auto_in_e_valid,
  input         auto_in_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [2:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [2:0]  auto_out_c_bits_size,
  output [6:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [2:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output        auto_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_bits_sink; // @[Nodes.scala 24:25]
  wire [32:0] _a_notFIFO_T_1 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T = auto_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_1 = {1'b0,$signed(_a_id_T)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_3 = $signed(_a_id_T_1) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_4 = $signed(_a_id_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _a_id_T_5 = auto_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_6 = {1'b0,$signed(_a_id_T_5)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_8 = $signed(_a_id_T_6) & 33'she0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_9 = $signed(_a_id_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _a_id_T_10 = auto_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_11 = {1'b0,$signed(_a_id_T_10)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_13 = $signed(_a_id_T_11) & 33'shc0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_14 = $signed(_a_id_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _a_id_T_15 = auto_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_16 = {1'b0,$signed(_a_id_T_15)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_18 = $signed(_a_id_T_16) & 33'shc0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_19 = $signed(_a_id_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _a_id_T_20 = auto_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _a_id_T_21 = {1'b0,$signed(_a_id_T_20)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_23 = $signed(_a_id_T_21) & 33'she0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_24 = $signed(_a_id_T_23) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _a_id_T_28 = _a_id_T_4 | _a_id_T_9 | _a_id_T_14 | _a_id_T_19 | _a_id_T_24; // @[Parameters.scala 615:89]
  wire [32:0] _a_id_T_32 = $signed(_a_notFIFO_T_1) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_33 = $signed(_a_id_T_32) == 33'sh0; // @[Parameters.scala 137:67]
  wire [1:0] _a_id_T_35 = _a_id_T_33 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_523 = {{1'd0}, _a_id_T_28}; // @[Mux.scala 27:72]
  wire [1:0] a_id = _GEN_523 | _a_id_T_35; // @[Mux.scala 27:72]
  wire  a_noDomain = a_id == 2'h0; // @[FIFOFixer.scala 55:29]
  wire  stalls_a_sel = auto_in_a_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg  flight_16; // @[FIFOFixer.scala 71:27]
  reg  flight_17; // @[FIFOFixer.scala 71:27]
  reg  flight_18; // @[FIFOFixer.scala 71:27]
  reg  flight_19; // @[FIFOFixer.scala 71:27]
  reg  flight_20; // @[FIFOFixer.scala 71:27]
  reg  flight_21; // @[FIFOFixer.scala 71:27]
  reg  flight_22; // @[FIFOFixer.scala 71:27]
  reg  flight_23; // @[FIFOFixer.scala 71:27]
  reg  flight_24; // @[FIFOFixer.scala 71:27]
  reg  flight_25; // @[FIFOFixer.scala 71:27]
  reg  flight_26; // @[FIFOFixer.scala 71:27]
  reg  flight_27; // @[FIFOFixer.scala 71:27]
  reg  flight_28; // @[FIFOFixer.scala 71:27]
  reg  flight_29; // @[FIFOFixer.scala 71:27]
  reg  flight_30; // @[FIFOFixer.scala 71:27]
  reg  flight_31; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id; // @[Reg.scala 15:16]
  wire  stalls_0 = stalls_a_sel & a_first & (flight_16 | flight_17 | flight_18 | flight_19 | flight_20 | flight_21 |
    flight_22 | flight_23 | flight_24 | flight_25 | flight_26 | flight_27 | flight_28 | flight_29 | flight_30 |
    flight_31) & (a_noDomain | stalls_id != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_1 = auto_in_a_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  reg  flight_32; // @[FIFOFixer.scala 71:27]
  reg  flight_33; // @[FIFOFixer.scala 71:27]
  reg  flight_34; // @[FIFOFixer.scala 71:27]
  reg  flight_35; // @[FIFOFixer.scala 71:27]
  reg  flight_36; // @[FIFOFixer.scala 71:27]
  reg  flight_37; // @[FIFOFixer.scala 71:27]
  reg  flight_38; // @[FIFOFixer.scala 71:27]
  reg  flight_39; // @[FIFOFixer.scala 71:27]
  reg  flight_40; // @[FIFOFixer.scala 71:27]
  reg  flight_41; // @[FIFOFixer.scala 71:27]
  reg  flight_42; // @[FIFOFixer.scala 71:27]
  reg  flight_43; // @[FIFOFixer.scala 71:27]
  reg  flight_44; // @[FIFOFixer.scala 71:27]
  reg  flight_45; // @[FIFOFixer.scala 71:27]
  reg  flight_46; // @[FIFOFixer.scala 71:27]
  reg  flight_47; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id_1; // @[Reg.scala 15:16]
  wire  stalls_1 = stalls_a_sel_1 & a_first & (flight_32 | flight_33 | flight_34 | flight_35 | flight_36 | flight_37 |
    flight_38 | flight_39 | flight_40 | flight_41 | flight_42 | flight_43 | flight_44 | flight_45 | flight_46 |
    flight_47) & (a_noDomain | stalls_id_1 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_2 = auto_in_a_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  reg  flight_48; // @[FIFOFixer.scala 71:27]
  reg  flight_49; // @[FIFOFixer.scala 71:27]
  reg  flight_50; // @[FIFOFixer.scala 71:27]
  reg  flight_51; // @[FIFOFixer.scala 71:27]
  reg  flight_52; // @[FIFOFixer.scala 71:27]
  reg  flight_53; // @[FIFOFixer.scala 71:27]
  reg  flight_54; // @[FIFOFixer.scala 71:27]
  reg  flight_55; // @[FIFOFixer.scala 71:27]
  reg  flight_56; // @[FIFOFixer.scala 71:27]
  reg  flight_57; // @[FIFOFixer.scala 71:27]
  reg  flight_58; // @[FIFOFixer.scala 71:27]
  reg  flight_59; // @[FIFOFixer.scala 71:27]
  reg  flight_60; // @[FIFOFixer.scala 71:27]
  reg  flight_61; // @[FIFOFixer.scala 71:27]
  reg  flight_62; // @[FIFOFixer.scala 71:27]
  reg  flight_63; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id_2; // @[Reg.scala 15:16]
  wire  stalls_2 = stalls_a_sel_2 & a_first & (flight_48 | flight_49 | flight_50 | flight_51 | flight_52 | flight_53 |
    flight_54 | flight_55 | flight_56 | flight_57 | flight_58 | flight_59 | flight_60 | flight_61 | flight_62 |
    flight_63) & (a_noDomain | stalls_id_2 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_3 = auto_in_a_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  reg  flight_64; // @[FIFOFixer.scala 71:27]
  reg  flight_65; // @[FIFOFixer.scala 71:27]
  reg  flight_66; // @[FIFOFixer.scala 71:27]
  reg  flight_67; // @[FIFOFixer.scala 71:27]
  reg  flight_68; // @[FIFOFixer.scala 71:27]
  reg  flight_69; // @[FIFOFixer.scala 71:27]
  reg  flight_70; // @[FIFOFixer.scala 71:27]
  reg  flight_71; // @[FIFOFixer.scala 71:27]
  reg  flight_72; // @[FIFOFixer.scala 71:27]
  reg  flight_73; // @[FIFOFixer.scala 71:27]
  reg  flight_74; // @[FIFOFixer.scala 71:27]
  reg  flight_75; // @[FIFOFixer.scala 71:27]
  reg  flight_76; // @[FIFOFixer.scala 71:27]
  reg  flight_77; // @[FIFOFixer.scala 71:27]
  reg  flight_78; // @[FIFOFixer.scala 71:27]
  reg  flight_79; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id_3; // @[Reg.scala 15:16]
  wire  stalls_3 = stalls_a_sel_3 & a_first & (flight_64 | flight_65 | flight_66 | flight_67 | flight_68 | flight_69 |
    flight_70 | flight_71 | flight_72 | flight_73 | flight_74 | flight_75 | flight_76 | flight_77 | flight_78 |
    flight_79) & (a_noDomain | stalls_id_3 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_4 = auto_in_a_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  reg  flight_80; // @[FIFOFixer.scala 71:27]
  reg  flight_81; // @[FIFOFixer.scala 71:27]
  reg  flight_82; // @[FIFOFixer.scala 71:27]
  reg  flight_83; // @[FIFOFixer.scala 71:27]
  reg  flight_84; // @[FIFOFixer.scala 71:27]
  reg  flight_85; // @[FIFOFixer.scala 71:27]
  reg  flight_86; // @[FIFOFixer.scala 71:27]
  reg  flight_87; // @[FIFOFixer.scala 71:27]
  reg  flight_88; // @[FIFOFixer.scala 71:27]
  reg  flight_89; // @[FIFOFixer.scala 71:27]
  reg  flight_90; // @[FIFOFixer.scala 71:27]
  reg  flight_91; // @[FIFOFixer.scala 71:27]
  reg  flight_92; // @[FIFOFixer.scala 71:27]
  reg  flight_93; // @[FIFOFixer.scala 71:27]
  reg  flight_94; // @[FIFOFixer.scala 71:27]
  reg  flight_95; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id_4; // @[Reg.scala 15:16]
  wire  stalls_4 = stalls_a_sel_4 & a_first & (flight_80 | flight_81 | flight_82 | flight_83 | flight_84 | flight_85 |
    flight_86 | flight_87 | flight_88 | flight_89 | flight_90 | flight_91 | flight_92 | flight_93 | flight_94 |
    flight_95) & (a_noDomain | stalls_id_4 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_5 = auto_in_a_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  reg  flight_96; // @[FIFOFixer.scala 71:27]
  reg  flight_97; // @[FIFOFixer.scala 71:27]
  reg  flight_98; // @[FIFOFixer.scala 71:27]
  reg  flight_99; // @[FIFOFixer.scala 71:27]
  reg  flight_100; // @[FIFOFixer.scala 71:27]
  reg  flight_101; // @[FIFOFixer.scala 71:27]
  reg  flight_102; // @[FIFOFixer.scala 71:27]
  reg  flight_103; // @[FIFOFixer.scala 71:27]
  reg  flight_104; // @[FIFOFixer.scala 71:27]
  reg  flight_105; // @[FIFOFixer.scala 71:27]
  reg  flight_106; // @[FIFOFixer.scala 71:27]
  reg  flight_107; // @[FIFOFixer.scala 71:27]
  reg  flight_108; // @[FIFOFixer.scala 71:27]
  reg  flight_109; // @[FIFOFixer.scala 71:27]
  reg  flight_110; // @[FIFOFixer.scala 71:27]
  reg  flight_111; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id_5; // @[Reg.scala 15:16]
  wire  stalls_5 = stalls_a_sel_5 & a_first & (flight_96 | flight_97 | flight_98 | flight_99 | flight_100 | flight_101
     | flight_102 | flight_103 | flight_104 | flight_105 | flight_106 | flight_107 | flight_108 | flight_109 |
    flight_110 | flight_111) & (a_noDomain | stalls_id_5 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_6 = auto_in_a_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  reg  flight_112; // @[FIFOFixer.scala 71:27]
  reg  flight_113; // @[FIFOFixer.scala 71:27]
  reg  flight_114; // @[FIFOFixer.scala 71:27]
  reg  flight_115; // @[FIFOFixer.scala 71:27]
  reg  flight_116; // @[FIFOFixer.scala 71:27]
  reg  flight_117; // @[FIFOFixer.scala 71:27]
  reg  flight_118; // @[FIFOFixer.scala 71:27]
  reg  flight_119; // @[FIFOFixer.scala 71:27]
  reg  flight_120; // @[FIFOFixer.scala 71:27]
  reg  flight_121; // @[FIFOFixer.scala 71:27]
  reg  flight_122; // @[FIFOFixer.scala 71:27]
  reg  flight_123; // @[FIFOFixer.scala 71:27]
  reg  flight_124; // @[FIFOFixer.scala 71:27]
  reg  flight_125; // @[FIFOFixer.scala 71:27]
  reg  flight_126; // @[FIFOFixer.scala 71:27]
  reg  flight_127; // @[FIFOFixer.scala 71:27]
  reg [1:0] stalls_id_6; // @[Reg.scala 15:16]
  wire  stalls_6 = stalls_a_sel_6 & a_first & (flight_112 | flight_113 | flight_114 | flight_115 | flight_116 |
    flight_117 | flight_118 | flight_119 | flight_120 | flight_121 | flight_122 | flight_123 | flight_124 | flight_125
     | flight_126 | flight_127) & (a_noDomain | stalls_id_6 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stall = stalls_0 | stalls_1 | stalls_2 | stalls_3 | stalls_4 | stalls_5 | stalls_6; // @[FIFOFixer.scala 83:49]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[FIFOFixer.scala 88:50]
  wire  bundleIn_0_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  wire  _a_first_T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _a_first_beats1_decode_T_1 = 13'h3f << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _a_first_beats1_decode_T_3 = ~_a_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] a_first_beats1_decode = _a_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  _d_first_T = auto_in_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  wire  d_first = d_first_first & auto_out_d_bits_opcode != 3'h6; // @[FIFOFixer.scala 67:42]
  wire  _GEN_146 = a_first & _a_first_T ? 7'h10 == auto_in_a_bits_source | flight_16 : flight_16; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_147 = a_first & _a_first_T ? 7'h11 == auto_in_a_bits_source | flight_17 : flight_17; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_148 = a_first & _a_first_T ? 7'h12 == auto_in_a_bits_source | flight_18 : flight_18; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_149 = a_first & _a_first_T ? 7'h13 == auto_in_a_bits_source | flight_19 : flight_19; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_150 = a_first & _a_first_T ? 7'h14 == auto_in_a_bits_source | flight_20 : flight_20; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_151 = a_first & _a_first_T ? 7'h15 == auto_in_a_bits_source | flight_21 : flight_21; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_152 = a_first & _a_first_T ? 7'h16 == auto_in_a_bits_source | flight_22 : flight_22; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_153 = a_first & _a_first_T ? 7'h17 == auto_in_a_bits_source | flight_23 : flight_23; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_154 = a_first & _a_first_T ? 7'h18 == auto_in_a_bits_source | flight_24 : flight_24; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_155 = a_first & _a_first_T ? 7'h19 == auto_in_a_bits_source | flight_25 : flight_25; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_156 = a_first & _a_first_T ? 7'h1a == auto_in_a_bits_source | flight_26 : flight_26; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_157 = a_first & _a_first_T ? 7'h1b == auto_in_a_bits_source | flight_27 : flight_27; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_158 = a_first & _a_first_T ? 7'h1c == auto_in_a_bits_source | flight_28 : flight_28; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_159 = a_first & _a_first_T ? 7'h1d == auto_in_a_bits_source | flight_29 : flight_29; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_160 = a_first & _a_first_T ? 7'h1e == auto_in_a_bits_source | flight_30 : flight_30; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_161 = a_first & _a_first_T ? 7'h1f == auto_in_a_bits_source | flight_31 : flight_31; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_162 = a_first & _a_first_T ? 7'h20 == auto_in_a_bits_source | flight_32 : flight_32; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_163 = a_first & _a_first_T ? 7'h21 == auto_in_a_bits_source | flight_33 : flight_33; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_164 = a_first & _a_first_T ? 7'h22 == auto_in_a_bits_source | flight_34 : flight_34; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_165 = a_first & _a_first_T ? 7'h23 == auto_in_a_bits_source | flight_35 : flight_35; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_166 = a_first & _a_first_T ? 7'h24 == auto_in_a_bits_source | flight_36 : flight_36; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_167 = a_first & _a_first_T ? 7'h25 == auto_in_a_bits_source | flight_37 : flight_37; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_168 = a_first & _a_first_T ? 7'h26 == auto_in_a_bits_source | flight_38 : flight_38; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_169 = a_first & _a_first_T ? 7'h27 == auto_in_a_bits_source | flight_39 : flight_39; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_170 = a_first & _a_first_T ? 7'h28 == auto_in_a_bits_source | flight_40 : flight_40; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_171 = a_first & _a_first_T ? 7'h29 == auto_in_a_bits_source | flight_41 : flight_41; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_172 = a_first & _a_first_T ? 7'h2a == auto_in_a_bits_source | flight_42 : flight_42; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_173 = a_first & _a_first_T ? 7'h2b == auto_in_a_bits_source | flight_43 : flight_43; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_174 = a_first & _a_first_T ? 7'h2c == auto_in_a_bits_source | flight_44 : flight_44; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_175 = a_first & _a_first_T ? 7'h2d == auto_in_a_bits_source | flight_45 : flight_45; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_176 = a_first & _a_first_T ? 7'h2e == auto_in_a_bits_source | flight_46 : flight_46; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_177 = a_first & _a_first_T ? 7'h2f == auto_in_a_bits_source | flight_47 : flight_47; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_178 = a_first & _a_first_T ? 7'h30 == auto_in_a_bits_source | flight_48 : flight_48; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_179 = a_first & _a_first_T ? 7'h31 == auto_in_a_bits_source | flight_49 : flight_49; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_180 = a_first & _a_first_T ? 7'h32 == auto_in_a_bits_source | flight_50 : flight_50; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_181 = a_first & _a_first_T ? 7'h33 == auto_in_a_bits_source | flight_51 : flight_51; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_182 = a_first & _a_first_T ? 7'h34 == auto_in_a_bits_source | flight_52 : flight_52; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_183 = a_first & _a_first_T ? 7'h35 == auto_in_a_bits_source | flight_53 : flight_53; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_184 = a_first & _a_first_T ? 7'h36 == auto_in_a_bits_source | flight_54 : flight_54; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_185 = a_first & _a_first_T ? 7'h37 == auto_in_a_bits_source | flight_55 : flight_55; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_186 = a_first & _a_first_T ? 7'h38 == auto_in_a_bits_source | flight_56 : flight_56; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_187 = a_first & _a_first_T ? 7'h39 == auto_in_a_bits_source | flight_57 : flight_57; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_188 = a_first & _a_first_T ? 7'h3a == auto_in_a_bits_source | flight_58 : flight_58; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_189 = a_first & _a_first_T ? 7'h3b == auto_in_a_bits_source | flight_59 : flight_59; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_190 = a_first & _a_first_T ? 7'h3c == auto_in_a_bits_source | flight_60 : flight_60; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_191 = a_first & _a_first_T ? 7'h3d == auto_in_a_bits_source | flight_61 : flight_61; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_192 = a_first & _a_first_T ? 7'h3e == auto_in_a_bits_source | flight_62 : flight_62; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_193 = a_first & _a_first_T ? 7'h3f == auto_in_a_bits_source | flight_63 : flight_63; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_194 = a_first & _a_first_T ? 7'h40 == auto_in_a_bits_source | flight_64 : flight_64; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_195 = a_first & _a_first_T ? 7'h41 == auto_in_a_bits_source | flight_65 : flight_65; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_196 = a_first & _a_first_T ? 7'h42 == auto_in_a_bits_source | flight_66 : flight_66; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_197 = a_first & _a_first_T ? 7'h43 == auto_in_a_bits_source | flight_67 : flight_67; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_198 = a_first & _a_first_T ? 7'h44 == auto_in_a_bits_source | flight_68 : flight_68; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_199 = a_first & _a_first_T ? 7'h45 == auto_in_a_bits_source | flight_69 : flight_69; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_200 = a_first & _a_first_T ? 7'h46 == auto_in_a_bits_source | flight_70 : flight_70; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_201 = a_first & _a_first_T ? 7'h47 == auto_in_a_bits_source | flight_71 : flight_71; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_202 = a_first & _a_first_T ? 7'h48 == auto_in_a_bits_source | flight_72 : flight_72; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_203 = a_first & _a_first_T ? 7'h49 == auto_in_a_bits_source | flight_73 : flight_73; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_204 = a_first & _a_first_T ? 7'h4a == auto_in_a_bits_source | flight_74 : flight_74; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_205 = a_first & _a_first_T ? 7'h4b == auto_in_a_bits_source | flight_75 : flight_75; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_206 = a_first & _a_first_T ? 7'h4c == auto_in_a_bits_source | flight_76 : flight_76; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_207 = a_first & _a_first_T ? 7'h4d == auto_in_a_bits_source | flight_77 : flight_77; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_208 = a_first & _a_first_T ? 7'h4e == auto_in_a_bits_source | flight_78 : flight_78; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_209 = a_first & _a_first_T ? 7'h4f == auto_in_a_bits_source | flight_79 : flight_79; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_210 = a_first & _a_first_T ? 7'h50 == auto_in_a_bits_source | flight_80 : flight_80; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_211 = a_first & _a_first_T ? 7'h51 == auto_in_a_bits_source | flight_81 : flight_81; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_212 = a_first & _a_first_T ? 7'h52 == auto_in_a_bits_source | flight_82 : flight_82; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_213 = a_first & _a_first_T ? 7'h53 == auto_in_a_bits_source | flight_83 : flight_83; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_214 = a_first & _a_first_T ? 7'h54 == auto_in_a_bits_source | flight_84 : flight_84; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_215 = a_first & _a_first_T ? 7'h55 == auto_in_a_bits_source | flight_85 : flight_85; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_216 = a_first & _a_first_T ? 7'h56 == auto_in_a_bits_source | flight_86 : flight_86; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_217 = a_first & _a_first_T ? 7'h57 == auto_in_a_bits_source | flight_87 : flight_87; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_218 = a_first & _a_first_T ? 7'h58 == auto_in_a_bits_source | flight_88 : flight_88; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_219 = a_first & _a_first_T ? 7'h59 == auto_in_a_bits_source | flight_89 : flight_89; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_220 = a_first & _a_first_T ? 7'h5a == auto_in_a_bits_source | flight_90 : flight_90; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_221 = a_first & _a_first_T ? 7'h5b == auto_in_a_bits_source | flight_91 : flight_91; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_222 = a_first & _a_first_T ? 7'h5c == auto_in_a_bits_source | flight_92 : flight_92; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_223 = a_first & _a_first_T ? 7'h5d == auto_in_a_bits_source | flight_93 : flight_93; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_224 = a_first & _a_first_T ? 7'h5e == auto_in_a_bits_source | flight_94 : flight_94; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_225 = a_first & _a_first_T ? 7'h5f == auto_in_a_bits_source | flight_95 : flight_95; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_226 = a_first & _a_first_T ? 7'h60 == auto_in_a_bits_source | flight_96 : flight_96; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_227 = a_first & _a_first_T ? 7'h61 == auto_in_a_bits_source | flight_97 : flight_97; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_228 = a_first & _a_first_T ? 7'h62 == auto_in_a_bits_source | flight_98 : flight_98; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_229 = a_first & _a_first_T ? 7'h63 == auto_in_a_bits_source | flight_99 : flight_99; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_230 = a_first & _a_first_T ? 7'h64 == auto_in_a_bits_source | flight_100 : flight_100; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_231 = a_first & _a_first_T ? 7'h65 == auto_in_a_bits_source | flight_101 : flight_101; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_232 = a_first & _a_first_T ? 7'h66 == auto_in_a_bits_source | flight_102 : flight_102; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_233 = a_first & _a_first_T ? 7'h67 == auto_in_a_bits_source | flight_103 : flight_103; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_234 = a_first & _a_first_T ? 7'h68 == auto_in_a_bits_source | flight_104 : flight_104; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_235 = a_first & _a_first_T ? 7'h69 == auto_in_a_bits_source | flight_105 : flight_105; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_236 = a_first & _a_first_T ? 7'h6a == auto_in_a_bits_source | flight_106 : flight_106; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_237 = a_first & _a_first_T ? 7'h6b == auto_in_a_bits_source | flight_107 : flight_107; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_238 = a_first & _a_first_T ? 7'h6c == auto_in_a_bits_source | flight_108 : flight_108; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_239 = a_first & _a_first_T ? 7'h6d == auto_in_a_bits_source | flight_109 : flight_109; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_240 = a_first & _a_first_T ? 7'h6e == auto_in_a_bits_source | flight_110 : flight_110; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_241 = a_first & _a_first_T ? 7'h6f == auto_in_a_bits_source | flight_111 : flight_111; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_242 = a_first & _a_first_T ? 7'h70 == auto_in_a_bits_source | flight_112 : flight_112; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_243 = a_first & _a_first_T ? 7'h71 == auto_in_a_bits_source | flight_113 : flight_113; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_244 = a_first & _a_first_T ? 7'h72 == auto_in_a_bits_source | flight_114 : flight_114; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_245 = a_first & _a_first_T ? 7'h73 == auto_in_a_bits_source | flight_115 : flight_115; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_246 = a_first & _a_first_T ? 7'h74 == auto_in_a_bits_source | flight_116 : flight_116; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_247 = a_first & _a_first_T ? 7'h75 == auto_in_a_bits_source | flight_117 : flight_117; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_248 = a_first & _a_first_T ? 7'h76 == auto_in_a_bits_source | flight_118 : flight_118; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_249 = a_first & _a_first_T ? 7'h77 == auto_in_a_bits_source | flight_119 : flight_119; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_250 = a_first & _a_first_T ? 7'h78 == auto_in_a_bits_source | flight_120 : flight_120; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_251 = a_first & _a_first_T ? 7'h79 == auto_in_a_bits_source | flight_121 : flight_121; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_252 = a_first & _a_first_T ? 7'h7a == auto_in_a_bits_source | flight_122 : flight_122; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_253 = a_first & _a_first_T ? 7'h7b == auto_in_a_bits_source | flight_123 : flight_123; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_254 = a_first & _a_first_T ? 7'h7c == auto_in_a_bits_source | flight_124 : flight_124; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_255 = a_first & _a_first_T ? 7'h7d == auto_in_a_bits_source | flight_125 : flight_125; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_256 = a_first & _a_first_T ? 7'h7e == auto_in_a_bits_source | flight_126 : flight_126; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _GEN_257 = a_first & _a_first_T ? 7'h7f == auto_in_a_bits_source | flight_127 : flight_127; // @[FIFOFixer.scala 72:37 FIFOFixer.scala 71:27]
  wire  _stalls_id_T_1 = _a_first_T & stalls_a_sel; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_5 = _a_first_T & stalls_a_sel_1; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_9 = _a_first_T & stalls_a_sel_2; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_13 = _a_first_T & stalls_a_sel_3; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_17 = _a_first_T & stalls_a_sel_4; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_21 = _a_first_T & stalls_a_sel_5; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_25 = _a_first_T & stalls_a_sel_6; // @[FIFOFixer.scala 77:49]
  TLMonitor_13 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_c_ready(monitor_io_in_c_ready),
    .io_in_c_valid(monitor_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_io_in_c_bits_address),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),
    .io_in_e_ready(monitor_io_in_e_ready),
    .io_in_e_valid(monitor_io_in_e_valid),
    .io_in_e_bits_sink(monitor_io_in_e_bits_sink)
  );
  assign auto_in_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  assign auto_in_c_ready = auto_out_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_e_ready = auto_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid & _bundleIn_0_a_ready_T; // @[FIFOFixer.scala 87:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_ready = auto_out_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_e_ready = auto_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_16 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h10 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_16 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_16 <= _GEN_146;
      end
    end else begin
      flight_16 <= _GEN_146;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_17 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h11 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_17 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_17 <= _GEN_147;
      end
    end else begin
      flight_17 <= _GEN_147;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_18 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h12 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_18 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_18 <= _GEN_148;
      end
    end else begin
      flight_18 <= _GEN_148;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_19 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h13 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_19 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_19 <= _GEN_149;
      end
    end else begin
      flight_19 <= _GEN_149;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_20 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h14 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_20 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_20 <= _GEN_150;
      end
    end else begin
      flight_20 <= _GEN_150;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_21 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h15 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_21 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_21 <= _GEN_151;
      end
    end else begin
      flight_21 <= _GEN_151;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_22 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h16 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_22 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_22 <= _GEN_152;
      end
    end else begin
      flight_22 <= _GEN_152;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_23 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h17 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_23 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_23 <= _GEN_153;
      end
    end else begin
      flight_23 <= _GEN_153;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_24 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h18 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_24 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_24 <= _GEN_154;
      end
    end else begin
      flight_24 <= _GEN_154;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_25 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h19 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_25 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_25 <= _GEN_155;
      end
    end else begin
      flight_25 <= _GEN_155;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_26 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h1a == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_26 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_26 <= _GEN_156;
      end
    end else begin
      flight_26 <= _GEN_156;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_27 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h1b == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_27 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_27 <= _GEN_157;
      end
    end else begin
      flight_27 <= _GEN_157;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_28 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h1c == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_28 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_28 <= _GEN_158;
      end
    end else begin
      flight_28 <= _GEN_158;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_29 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h1d == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_29 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_29 <= _GEN_159;
      end
    end else begin
      flight_29 <= _GEN_159;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_30 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h1e == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_30 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_30 <= _GEN_160;
      end
    end else begin
      flight_30 <= _GEN_160;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_31 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h1f == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_31 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_31 <= _GEN_161;
      end
    end else begin
      flight_31 <= _GEN_161;
    end
    if (_stalls_id_T_1) begin // @[Reg.scala 16:19]
      stalls_id <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_32 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h20 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_32 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_32 <= _GEN_162;
      end
    end else begin
      flight_32 <= _GEN_162;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_33 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h21 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_33 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_33 <= _GEN_163;
      end
    end else begin
      flight_33 <= _GEN_163;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_34 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h22 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_34 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_34 <= _GEN_164;
      end
    end else begin
      flight_34 <= _GEN_164;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_35 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h23 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_35 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_35 <= _GEN_165;
      end
    end else begin
      flight_35 <= _GEN_165;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_36 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h24 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_36 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_36 <= _GEN_166;
      end
    end else begin
      flight_36 <= _GEN_166;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_37 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h25 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_37 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_37 <= _GEN_167;
      end
    end else begin
      flight_37 <= _GEN_167;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_38 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h26 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_38 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_38 <= _GEN_168;
      end
    end else begin
      flight_38 <= _GEN_168;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_39 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h27 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_39 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_39 <= _GEN_169;
      end
    end else begin
      flight_39 <= _GEN_169;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_40 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h28 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_40 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_40 <= _GEN_170;
      end
    end else begin
      flight_40 <= _GEN_170;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_41 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h29 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_41 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_41 <= _GEN_171;
      end
    end else begin
      flight_41 <= _GEN_171;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_42 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h2a == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_42 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_42 <= _GEN_172;
      end
    end else begin
      flight_42 <= _GEN_172;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_43 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h2b == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_43 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_43 <= _GEN_173;
      end
    end else begin
      flight_43 <= _GEN_173;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_44 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h2c == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_44 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_44 <= _GEN_174;
      end
    end else begin
      flight_44 <= _GEN_174;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_45 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h2d == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_45 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_45 <= _GEN_175;
      end
    end else begin
      flight_45 <= _GEN_175;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_46 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h2e == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_46 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_46 <= _GEN_176;
      end
    end else begin
      flight_46 <= _GEN_176;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_47 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h2f == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_47 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_47 <= _GEN_177;
      end
    end else begin
      flight_47 <= _GEN_177;
    end
    if (_stalls_id_T_5) begin // @[Reg.scala 16:19]
      stalls_id_1 <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_48 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h30 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_48 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_48 <= _GEN_178;
      end
    end else begin
      flight_48 <= _GEN_178;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_49 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h31 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_49 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_49 <= _GEN_179;
      end
    end else begin
      flight_49 <= _GEN_179;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_50 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h32 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_50 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_50 <= _GEN_180;
      end
    end else begin
      flight_50 <= _GEN_180;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_51 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h33 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_51 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_51 <= _GEN_181;
      end
    end else begin
      flight_51 <= _GEN_181;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_52 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h34 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_52 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_52 <= _GEN_182;
      end
    end else begin
      flight_52 <= _GEN_182;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_53 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h35 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_53 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_53 <= _GEN_183;
      end
    end else begin
      flight_53 <= _GEN_183;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_54 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h36 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_54 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_54 <= _GEN_184;
      end
    end else begin
      flight_54 <= _GEN_184;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_55 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h37 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_55 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_55 <= _GEN_185;
      end
    end else begin
      flight_55 <= _GEN_185;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_56 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h38 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_56 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_56 <= _GEN_186;
      end
    end else begin
      flight_56 <= _GEN_186;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_57 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h39 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_57 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_57 <= _GEN_187;
      end
    end else begin
      flight_57 <= _GEN_187;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_58 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h3a == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_58 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_58 <= _GEN_188;
      end
    end else begin
      flight_58 <= _GEN_188;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_59 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h3b == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_59 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_59 <= _GEN_189;
      end
    end else begin
      flight_59 <= _GEN_189;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_60 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h3c == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_60 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_60 <= _GEN_190;
      end
    end else begin
      flight_60 <= _GEN_190;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_61 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h3d == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_61 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_61 <= _GEN_191;
      end
    end else begin
      flight_61 <= _GEN_191;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_62 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h3e == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_62 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_62 <= _GEN_192;
      end
    end else begin
      flight_62 <= _GEN_192;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_63 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h3f == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_63 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_63 <= _GEN_193;
      end
    end else begin
      flight_63 <= _GEN_193;
    end
    if (_stalls_id_T_9) begin // @[Reg.scala 16:19]
      stalls_id_2 <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_64 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h40 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_64 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_64 <= _GEN_194;
      end
    end else begin
      flight_64 <= _GEN_194;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_65 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h41 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_65 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_65 <= _GEN_195;
      end
    end else begin
      flight_65 <= _GEN_195;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_66 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h42 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_66 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_66 <= _GEN_196;
      end
    end else begin
      flight_66 <= _GEN_196;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_67 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h43 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_67 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_67 <= _GEN_197;
      end
    end else begin
      flight_67 <= _GEN_197;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_68 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h44 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_68 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_68 <= _GEN_198;
      end
    end else begin
      flight_68 <= _GEN_198;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_69 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h45 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_69 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_69 <= _GEN_199;
      end
    end else begin
      flight_69 <= _GEN_199;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_70 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h46 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_70 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_70 <= _GEN_200;
      end
    end else begin
      flight_70 <= _GEN_200;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_71 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h47 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_71 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_71 <= _GEN_201;
      end
    end else begin
      flight_71 <= _GEN_201;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_72 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h48 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_72 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_72 <= _GEN_202;
      end
    end else begin
      flight_72 <= _GEN_202;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_73 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h49 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_73 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_73 <= _GEN_203;
      end
    end else begin
      flight_73 <= _GEN_203;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_74 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h4a == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_74 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_74 <= _GEN_204;
      end
    end else begin
      flight_74 <= _GEN_204;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_75 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h4b == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_75 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_75 <= _GEN_205;
      end
    end else begin
      flight_75 <= _GEN_205;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_76 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h4c == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_76 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_76 <= _GEN_206;
      end
    end else begin
      flight_76 <= _GEN_206;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_77 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h4d == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_77 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_77 <= _GEN_207;
      end
    end else begin
      flight_77 <= _GEN_207;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_78 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h4e == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_78 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_78 <= _GEN_208;
      end
    end else begin
      flight_78 <= _GEN_208;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_79 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h4f == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_79 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_79 <= _GEN_209;
      end
    end else begin
      flight_79 <= _GEN_209;
    end
    if (_stalls_id_T_13) begin // @[Reg.scala 16:19]
      stalls_id_3 <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_80 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h50 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_80 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_80 <= _GEN_210;
      end
    end else begin
      flight_80 <= _GEN_210;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_81 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h51 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_81 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_81 <= _GEN_211;
      end
    end else begin
      flight_81 <= _GEN_211;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_82 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h52 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_82 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_82 <= _GEN_212;
      end
    end else begin
      flight_82 <= _GEN_212;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_83 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h53 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_83 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_83 <= _GEN_213;
      end
    end else begin
      flight_83 <= _GEN_213;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_84 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h54 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_84 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_84 <= _GEN_214;
      end
    end else begin
      flight_84 <= _GEN_214;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_85 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h55 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_85 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_85 <= _GEN_215;
      end
    end else begin
      flight_85 <= _GEN_215;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_86 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h56 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_86 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_86 <= _GEN_216;
      end
    end else begin
      flight_86 <= _GEN_216;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_87 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h57 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_87 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_87 <= _GEN_217;
      end
    end else begin
      flight_87 <= _GEN_217;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_88 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h58 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_88 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_88 <= _GEN_218;
      end
    end else begin
      flight_88 <= _GEN_218;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_89 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h59 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_89 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_89 <= _GEN_219;
      end
    end else begin
      flight_89 <= _GEN_219;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_90 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h5a == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_90 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_90 <= _GEN_220;
      end
    end else begin
      flight_90 <= _GEN_220;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_91 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h5b == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_91 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_91 <= _GEN_221;
      end
    end else begin
      flight_91 <= _GEN_221;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_92 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h5c == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_92 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_92 <= _GEN_222;
      end
    end else begin
      flight_92 <= _GEN_222;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_93 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h5d == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_93 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_93 <= _GEN_223;
      end
    end else begin
      flight_93 <= _GEN_223;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_94 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h5e == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_94 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_94 <= _GEN_224;
      end
    end else begin
      flight_94 <= _GEN_224;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_95 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h5f == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_95 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_95 <= _GEN_225;
      end
    end else begin
      flight_95 <= _GEN_225;
    end
    if (_stalls_id_T_17) begin // @[Reg.scala 16:19]
      stalls_id_4 <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_96 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h60 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_96 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_96 <= _GEN_226;
      end
    end else begin
      flight_96 <= _GEN_226;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_97 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h61 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_97 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_97 <= _GEN_227;
      end
    end else begin
      flight_97 <= _GEN_227;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_98 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h62 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_98 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_98 <= _GEN_228;
      end
    end else begin
      flight_98 <= _GEN_228;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_99 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h63 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_99 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_99 <= _GEN_229;
      end
    end else begin
      flight_99 <= _GEN_229;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_100 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h64 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_100 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_100 <= _GEN_230;
      end
    end else begin
      flight_100 <= _GEN_230;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_101 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h65 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_101 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_101 <= _GEN_231;
      end
    end else begin
      flight_101 <= _GEN_231;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_102 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h66 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_102 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_102 <= _GEN_232;
      end
    end else begin
      flight_102 <= _GEN_232;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_103 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h67 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_103 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_103 <= _GEN_233;
      end
    end else begin
      flight_103 <= _GEN_233;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_104 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h68 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_104 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_104 <= _GEN_234;
      end
    end else begin
      flight_104 <= _GEN_234;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_105 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h69 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_105 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_105 <= _GEN_235;
      end
    end else begin
      flight_105 <= _GEN_235;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_106 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h6a == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_106 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_106 <= _GEN_236;
      end
    end else begin
      flight_106 <= _GEN_236;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_107 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h6b == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_107 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_107 <= _GEN_237;
      end
    end else begin
      flight_107 <= _GEN_237;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_108 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h6c == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_108 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_108 <= _GEN_238;
      end
    end else begin
      flight_108 <= _GEN_238;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_109 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h6d == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_109 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_109 <= _GEN_239;
      end
    end else begin
      flight_109 <= _GEN_239;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_110 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h6e == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_110 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_110 <= _GEN_240;
      end
    end else begin
      flight_110 <= _GEN_240;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_111 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h6f == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_111 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_111 <= _GEN_241;
      end
    end else begin
      flight_111 <= _GEN_241;
    end
    if (_stalls_id_T_21) begin // @[Reg.scala 16:19]
      stalls_id_5 <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_112 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h70 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_112 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_112 <= _GEN_242;
      end
    end else begin
      flight_112 <= _GEN_242;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_113 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h71 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_113 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_113 <= _GEN_243;
      end
    end else begin
      flight_113 <= _GEN_243;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_114 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h72 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_114 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_114 <= _GEN_244;
      end
    end else begin
      flight_114 <= _GEN_244;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_115 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h73 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_115 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_115 <= _GEN_245;
      end
    end else begin
      flight_115 <= _GEN_245;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_116 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h74 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_116 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_116 <= _GEN_246;
      end
    end else begin
      flight_116 <= _GEN_246;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_117 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h75 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_117 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_117 <= _GEN_247;
      end
    end else begin
      flight_117 <= _GEN_247;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_118 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h76 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_118 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_118 <= _GEN_248;
      end
    end else begin
      flight_118 <= _GEN_248;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_119 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h77 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_119 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_119 <= _GEN_249;
      end
    end else begin
      flight_119 <= _GEN_249;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_120 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h78 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_120 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_120 <= _GEN_250;
      end
    end else begin
      flight_120 <= _GEN_250;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_121 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h79 == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_121 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_121 <= _GEN_251;
      end
    end else begin
      flight_121 <= _GEN_251;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_122 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h7a == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_122 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_122 <= _GEN_252;
      end
    end else begin
      flight_122 <= _GEN_252;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_123 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h7b == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_123 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_123 <= _GEN_253;
      end
    end else begin
      flight_123 <= _GEN_253;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_124 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h7c == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_124 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_124 <= _GEN_254;
      end
    end else begin
      flight_124 <= _GEN_254;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_125 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h7d == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_125 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_125 <= _GEN_255;
      end
    end else begin
      flight_125 <= _GEN_255;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_126 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h7e == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_126 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_126 <= _GEN_256;
      end
    end else begin
      flight_126 <= _GEN_256;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_127 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin // @[FIFOFixer.scala 73:37]
      if (7'h7f == auto_out_d_bits_source) begin // @[FIFOFixer.scala 73:64]
        flight_127 <= 1'h0; // @[FIFOFixer.scala 73:64]
      end else begin
        flight_127 <= _GEN_257;
      end
    end else begin
      flight_127 <= _GEN_257;
    end
    if (_stalls_id_T_25) begin // @[Reg.scala 16:19]
      stalls_id_6 <= a_id; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  flight_16 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  flight_17 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  flight_18 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  flight_19 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  flight_20 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  flight_21 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  flight_22 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  flight_23 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  flight_24 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  flight_25 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  flight_26 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  flight_27 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  flight_28 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  flight_29 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  flight_30 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  flight_31 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  stalls_id = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  flight_32 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  flight_33 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  flight_34 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  flight_35 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  flight_36 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  flight_37 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  flight_38 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  flight_39 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  flight_40 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  flight_41 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  flight_42 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  flight_43 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  flight_44 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  flight_45 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  flight_46 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  flight_47 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  stalls_id_1 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  flight_48 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  flight_49 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  flight_50 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  flight_51 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  flight_52 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  flight_53 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  flight_54 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  flight_55 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  flight_56 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  flight_57 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  flight_58 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  flight_59 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  flight_60 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  flight_61 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  flight_62 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  flight_63 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  stalls_id_2 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  flight_64 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  flight_65 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  flight_66 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  flight_67 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  flight_68 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  flight_69 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  flight_70 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  flight_71 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  flight_72 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  flight_73 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  flight_74 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  flight_75 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  flight_76 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  flight_77 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  flight_78 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  flight_79 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  stalls_id_3 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  flight_80 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  flight_81 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  flight_82 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  flight_83 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  flight_84 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  flight_85 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  flight_86 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  flight_87 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  flight_88 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  flight_89 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  flight_90 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  flight_91 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  flight_92 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  flight_93 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  flight_94 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  flight_95 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  stalls_id_4 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  flight_96 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  flight_97 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  flight_98 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  flight_99 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  flight_100 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  flight_101 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  flight_102 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  flight_103 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  flight_104 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  flight_105 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  flight_106 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  flight_107 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  flight_108 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  flight_109 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  flight_110 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  flight_111 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  stalls_id_5 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  flight_112 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  flight_113 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  flight_114 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  flight_115 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  flight_116 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  flight_117 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  flight_118 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  flight_119 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  flight_120 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  flight_121 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  flight_122 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  flight_123 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  flight_124 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  flight_125 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  flight_126 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  flight_127 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  stalls_id_6 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  d_first_counter = _RAND_120[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_14(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [5:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [2:0]  io_in_c_bits_size,
  input  [5:0]  io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [5:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input         io_in_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [255:0] _RAND_19;
  reg [255:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [255:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_86 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_2 = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_3 = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_4 = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_5 = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_lo = mask_acc_2 | mask_size_2 & mask_eq_6; // @[Misc.scala 214:29]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_hi = mask_acc_2 | mask_size_2 & mask_eq_7; // @[Misc.scala 214:29]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_lo = mask_acc_3 | mask_size_2 & mask_eq_8; // @[Misc.scala 214:29]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_hi = mask_acc_3 | mask_size_2 & mask_eq_9; // @[Misc.scala 214:29]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_lo = mask_acc_4 | mask_size_2 & mask_eq_10; // @[Misc.scala 214:29]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_hi = mask_acc_4 | mask_size_2 & mask_eq_11; // @[Misc.scala 214:29]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_lo = mask_acc_5 | mask_size_2 & mask_eq_12; // @[Misc.scala 214:29]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_hi = mask_acc_5 | mask_size_2 & mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire [31:0] _T_180 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_181 = {1'b0,$signed(_T_180)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_183 = $signed(_T_181) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_184 = $signed(_T_183) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_185 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_186 = {1'b0,$signed(_T_185)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_188 = $signed(_T_186) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_189 = $signed(_T_188) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_190 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_191 = {1'b0,$signed(_T_190)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_193 = $signed(_T_191) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_194 = $signed(_T_193) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_195 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_196 = {1'b0,$signed(_T_195)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_198 = $signed(_T_196) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_199 = $signed(_T_198) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_200 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_201 = {1'b0,$signed(_T_200)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_203 = $signed(_T_201) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_204 = $signed(_T_203) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_211 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_214 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_215 = {1'b0,$signed(_T_214)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_217 = $signed(_T_215) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_218 = $signed(_T_217) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_219 = _T_211 & _T_218; // @[Parameters.scala 670:56]
  wire  _T_222 = source_ok & _T_219; // @[Monitor.scala 82:72]
  wire  _T_277 = _source_ok_T_1 & _T_211; // @[Mux.scala 27:72]
  wire  _T_330 = _T_218 | _T_184 | _T_189 | _T_194 | _T_199 | _T_204; // @[Parameters.scala 671:42]
  wire  _T_333 = _T_277 & _T_330; // @[Monitor.scala 83:78]
  wire  _T_347 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [7:0] _T_351 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_352 = _T_351 == 8'h0; // @[Monitor.scala 88:31]
  wire  _T_360 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_593 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_606 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_709 = _T_211 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_720 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_724 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_732 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_834 = source_ok & _T_709; // @[Monitor.scala 115:71]
  wire  _T_852 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [7:0] _T_968 = ~mask; // @[Monitor.scala 127:33]
  wire [7:0] _T_969 = io_in_a_bits_mask & _T_968; // @[Monitor.scala 127:31]
  wire  _T_970 = _T_969 == 8'h0; // @[Monitor.scala 127:40]
  wire  _T_974 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_1036 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_1074 = _T_1036 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_1076 = source_ok & _T_1074; // @[Monitor.scala 131:74]
  wire  _T_1086 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_1094 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_1206 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_1214 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1326 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1338 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1342 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1346 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27]
  wire  _T_1350 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_1354 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1358 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1362 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1373 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_1377 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_1390 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1410 = _T_1358 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1419 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1436 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1454 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _source_ok_T_109 = io_in_c_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_115 = io_in_c_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_121 = io_in_c_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_127 = io_in_c_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_133 = io_in_c_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_139 = io_in_c_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_145 = io_in_c_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_151 = io_in_c_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_2 = _source_ok_T_109 | _source_ok_T_115 | _source_ok_T_121 | _source_ok_T_127 | _source_ok_T_133 |
    _source_ok_T_139 | _source_ok_T_145 | _source_ok_T_151; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_7 = 13'h3f << io_in_c_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask_2 = ~_is_aligned_mask_T_7[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_87 = {{26'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T_2 = io_in_c_bits_address & _GEN_87; // @[Edges.scala 20:16]
  wire  is_aligned_2 = _is_aligned_T_2 == 32'h0; // @[Edges.scala 20:24]
  wire [31:0] _address_ok_T_34 = io_in_c_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_35 = {1'b0,$signed(_address_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_37 = $signed(_address_ok_T_35) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_38 = $signed(_address_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_39 = io_in_c_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_40 = {1'b0,$signed(_address_ok_T_39)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_42 = $signed(_address_ok_T_40) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_43 = $signed(_address_ok_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_44 = io_in_c_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_45 = {1'b0,$signed(_address_ok_T_44)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_47 = $signed(_address_ok_T_45) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_48 = $signed(_address_ok_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_49 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_50 = {1'b0,$signed(_address_ok_T_49)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_52 = $signed(_address_ok_T_50) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_53 = $signed(_address_ok_T_52) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_54 = io_in_c_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_55 = {1'b0,$signed(_address_ok_T_54)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_57 = $signed(_address_ok_T_55) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_58 = $signed(_address_ok_T_57) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _address_ok_T_62 = _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 | _address_ok_T_58; // @[Parameters.scala 598:92]
  wire [31:0] _address_ok_T_63 = io_in_c_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_64 = {1'b0,$signed(_address_ok_T_63)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_66 = $signed(_address_ok_T_64) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_67 = $signed(_address_ok_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  wire  address_ok_1 = _address_ok_T_62 | _address_ok_T_67; // @[Parameters.scala 622:64]
  wire  _T_2224 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  wire  _T_2231 = io_in_c_bits_size >= 3'h3; // @[Monitor.scala 245:30]
  wire  _T_2238 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  wire  _T_2246 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  wire  _T_2264 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  wire  _T_2357 = io_in_c_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_2365 = _T_2357 & _address_ok_T_67; // @[Parameters.scala 670:56]
  wire  _T_2368 = source_ok_2 & _T_2365; // @[Monitor.scala 260:78]
  wire  _T_2423 = _source_ok_T_109 & _T_2357; // @[Mux.scala 27:72]
  wire  _T_2476 = _address_ok_T_67 | _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 |
    _address_ok_T_58; // @[Parameters.scala 671:42]
  wire  _T_2479 = _T_2423 & _T_2476; // @[Monitor.scala 261:78]
  wire  _T_2501 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  wire  _T_2734 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  wire  _T_2744 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  wire  _T_2752 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  wire  _T_2766 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  wire  sink_ok_1 = io_in_e_bits_sink < 1'h1; // @[Monitor.scala 364:31]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [5:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_2788 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_2789 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_2793 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_2797 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_2801 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_2805 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [5:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_2812 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_2813 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_2817 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_2821 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_2825 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_2833 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  wire  _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  wire [2:0] c_first_beats1_decode = is_aligned_mask_2[5:3]; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  reg [2:0] c_first_counter; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1 = c_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  c_first = c_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [2:0] size_3; // @[Monitor.scala 514:22]
  reg [5:0] source_3; // @[Monitor.scala 515:22]
  reg [31:0] address_2; // @[Monitor.scala 516:22]
  wire  _T_2864 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  wire  _T_2865 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  wire  _T_2869 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  wire  _T_2873 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  wire  _T_2877 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  wire  _T_2881 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  reg [63:0] inflight; // @[Monitor.scala 611:27]
  reg [255:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [255:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  wire [7:0] _GEN_88 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [8:0] _a_opcode_lookup_T = {{1'd0}, _GEN_88}; // @[Monitor.scala 634:69]
  wire [255:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [255:0] _GEN_89 = {{240'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [255:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_89; // @[Monitor.scala 634:97]
  wire [255:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[255:1]}; // @[Monitor.scala 634:152]
  wire [255:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [255:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 638:91]
  wire [255:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[255:1]}; // @[Monitor.scala 638:144]
  wire  _T_2887 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [63:0] _a_set_wo_ready_T = 64'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 64'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_2890 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [7:0] _GEN_94 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [8:0] _a_opcodes_set_T = {{1'd0}, _GEN_94}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [514:0] _GEN_95 = {{511'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [514:0] _a_opcodes_set_T_1 = _GEN_95 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [514:0] _GEN_97 = {{511'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [514:0] _a_sizes_set_T_1 = _GEN_97 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [63:0] _T_2892 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_2894 = ~_T_2892[0]; // @[Monitor.scala 658:17]
  wire [63:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 64'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [514:0] _GEN_31 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 515'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [514:0] _GEN_32 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 515'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_2898 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_2900 = ~_T_1342; // @[Monitor.scala 671:74]
  wire  _T_2901 = io_in_d_valid & d_first_1 & ~_T_1342; // @[Monitor.scala 671:71]
  wire [63:0] _d_clr_wo_ready_T = 64'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [526:0] _GEN_99 = {{511'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [526:0] _d_opcodes_clr_T_5 = _GEN_99 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [63:0] d_clr = _d_first_T & d_first_1 & _T_2900 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [526:0] _GEN_35 = _d_first_T & d_first_1 & _T_2900 ? _d_opcodes_clr_T_5 : 527'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_2887 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [63:0] _T_2911 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_2913 = _T_2911[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_2918 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_2919 = io_in_d_bits_opcode == _GEN_44 | _T_2918; // @[Monitor.scala 685:77]
  wire  _T_2923 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_2930 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_2931 = io_in_d_bits_opcode == _GEN_60 | _T_2930; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_102 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_2935 = _GEN_102 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_2945 = _T_2898 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_2900; // @[Monitor.scala 694:116]
  wire  _T_2946 = ~io_in_d_ready; // @[Monitor.scala 695:15]
  wire  _T_2947 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_2954 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [63:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [63:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [63:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [255:0] a_opcodes_set = _GEN_31[255:0];
  wire [255:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [255:0] d_opcodes_clr = _GEN_35[255:0];
  wire [255:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [255:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [255:0] a_sizes_set = _GEN_32[255:0];
  wire [255:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [255:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_2963 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [63:0] inflight_1; // @[Monitor.scala 723:35]
  reg [255:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [2:0] c_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1_1 = c_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  c_first_1 = c_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25]
  wire [255:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [255:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 747:93]
  wire [255:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[255:1]}; // @[Monitor.scala 747:146]
  wire  _T_2973 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  _T_2974 = io_in_c_valid & c_first_1 & _T_2973; // @[Monitor.scala 756:37]
  wire [63:0] _c_set_wo_ready_T = 64'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] c_set_wo_ready = io_in_c_valid & c_first_1 & _T_2973 ? _c_set_wo_ready_T : 64'h0; // @[Monitor.scala 756:71 Monitor.scala 757:22]
  wire  _T_2980 = _c_first_T & c_first_1 & _T_2973; // @[Monitor.scala 760:38]
  wire [3:0] _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  wire [3:0] _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 4'h1; // @[Monitor.scala 763:59]
  wire [7:0] _GEN_109 = {io_in_c_bits_source, 2'h0}; // @[Monitor.scala 764:79]
  wire [8:0] _c_opcodes_set_T = {{1'd0}, _GEN_109}; // @[Monitor.scala 764:79]
  wire [3:0] c_sizes_set_interm = _c_first_T & c_first_1 & _T_2973 ? _c_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 760:72 Monitor.scala 763:28]
  wire [514:0] _GEN_112 = {{511'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  wire [514:0] _c_sizes_set_T_1 = _GEN_112 << _c_opcodes_set_T; // @[Monitor.scala 765:52]
  wire [63:0] _T_2981 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  wire  _T_2983 = ~_T_2981[0]; // @[Monitor.scala 766:17]
  wire [63:0] c_set = _c_first_T & c_first_1 & _T_2973 ? _c_set_wo_ready_T : 64'h0; // @[Monitor.scala 760:72 Monitor.scala 761:28]
  wire [514:0] _GEN_77 = _c_first_T & c_first_1 & _T_2973 ? _c_sizes_set_T_1 : 515'h0; // @[Monitor.scala 760:72 Monitor.scala 765:28]
  wire  _T_2987 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  wire  _T_2989 = io_in_d_valid & d_first_2 & _T_1342; // @[Monitor.scala 779:71]
  wire [63:0] d_clr_wo_ready_1 = io_in_d_valid & d_first_2 & _T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 779:89 Monitor.scala 780:22]
  wire [63:0] d_clr_1 = _d_first_T & d_first_2 & _T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [526:0] _GEN_80 = _d_first_T & d_first_2 & _T_1342 ? _d_opcodes_clr_T_5 : 527'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire  _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1 = _T_2974 & io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:88]
  wire [63:0] _T_2997 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire  _T_2999 = _T_2997[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  wire  _T_3003 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_3007 = _GEN_102 == c_size_lookup; // @[Monitor.scala 795:36]
  wire  _T_3016 = _T_2987 & c_first_1 & io_in_c_valid & _same_cycle_resp_T_8 & _T_1342; // @[Monitor.scala 799:116]
  wire  _T_3018 = _T_2946 | io_in_c_ready; // @[Monitor.scala 800:32]
  wire  _T_3022 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  wire  _T_3023 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  wire [63:0] _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  wire [63:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [63:0] _inflight_T_5 = _inflight_T_3 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [255:0] d_opcodes_clr_1 = _GEN_80[255:0];
  wire [255:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [255:0] c_sizes_set = _GEN_77[255:0];
  wire [255:0] _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  wire [255:0] _inflight_sizes_T_5 = _inflight_sizes_T_3 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_3032 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [2:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_3 = d_first_counter_3 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 3'h0; // @[Edges.scala 230:25]
  wire  _T_3044 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_3045 = _d_first_T & d_first_3 & _T_3044; // @[Monitor.scala 829:38]
  wire  _T_3048 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = _d_first_T & d_first_3 & _T_3044 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  _T_3052 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _e_clr_T = 2'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  wire  d_set = _GEN_84[0];
  wire  _T_3056 = (d_set | inflight_2) >> io_in_e_bits_sink; // @[Monitor.scala 837:35]
  wire [1:0] _GEN_85 = _T_3052 ? _e_clr_T : 2'h0; // @[Monitor.scala 835:73 Monitor.scala 836:13]
  wire  e_clr = _GEN_85[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 3'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      opcode_3 <= io_in_c_bits_opcode; // @[Monitor.scala 525:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      param_3 <= io_in_c_bits_param; // @[Monitor.scala 526:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      size_3 <= io_in_c_bits_size; // @[Monitor.scala 527:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      source_3 <= io_in_c_bits_source; // @[Monitor.scala 528:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      address_2 <= io_in_c_bits_address; // @[Monitor.scala 529:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 64'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 256'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 256'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 64'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 256'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first_1) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 3'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_c_first_T | _d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= (inflight_2 | d_set) & ~e_clr; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 3'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1326 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1326 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1338 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1338 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1358 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1358 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1373 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1373 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1377 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1377 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1373 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1373 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1377 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1377 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1410 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1410 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2368 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2368 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2479 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2479 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid report param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2368 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2368 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2479 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2479 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channels carries invalid sink ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2789 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2789 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2793 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2793 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2797 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2797 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2801 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2805 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2813 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2813 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2817 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2817 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2821 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2821 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2825 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2825 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2833 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2833 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2865 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2865 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2869 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2869 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2873 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2873 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2877 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2877 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2881 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2881 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2890 & ~(_T_2894 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2890 & ~(_T_2894 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~(_T_2913 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~(_T_2913 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2919 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2919 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2923 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2923 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2931 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2931 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2935 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2935 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2945 & ~(_T_2947 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2945 & ~(_T_2947 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2954 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2954 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2963 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2963 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2980 & ~(_T_2983 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel re-used a source ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2980 & ~(_T_2983 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & ~(_T_2999 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & ~(_T_2999 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & same_cycle_resp_1 & ~(_T_3003 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & same_cycle_resp_1 & ~(_T_3003 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & ~same_cycle_resp_1 & ~(_T_3007 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & ~same_cycle_resp_1 & ~(_T_3007 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3016 & ~(_T_3018 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3016 & ~(_T_3018 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3022 & ~(_T_3023 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3022 & ~(_T_3023 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_3032 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_3032 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3045 & ~(_T_3048 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3045 & ~(_T_3048 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3052 & ~(_T_3056 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:98)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3052 & ~(_T_3056 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  c_first_counter = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  opcode_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  param_3 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  size_3 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  source_3 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  address_2 = _RAND_17[31:0];
  _RAND_18 = {2{`RANDOM}};
  inflight = _RAND_18[63:0];
  _RAND_19 = {8{`RANDOM}};
  inflight_opcodes = _RAND_19[255:0];
  _RAND_20 = {8{`RANDOM}};
  inflight_sizes = _RAND_20[255:0];
  _RAND_21 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  watchdog = _RAND_23[31:0];
  _RAND_24 = {2{`RANDOM}};
  inflight_1 = _RAND_24[63:0];
  _RAND_25 = {8{`RANDOM}};
  inflight_sizes_1 = _RAND_25[255:0];
  _RAND_26 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  watchdog_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inflight_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_30[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_1(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_size,
  input  [5:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_size,
  output [5:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [5:0] saved_source; // @[Repeater.scala 20:18]
  reg [31:0] saved_address; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 28:38 Repeater.scala 28:45 Repeater.scala 19:21]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign io_full = full; // @[Repeater.scala 26:11]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin // @[Repeater.scala 29:38]
      full <= 1'h0; // @[Repeater.scala 29:45]
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_size = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_source = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  saved_address = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLHintHandler(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [5:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [2:0]  auto_in_c_bits_size,
  input  [5:0]  auto_in_c_bits_source,
  input  [31:0] auto_in_c_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [5:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  output        auto_in_e_ready,
  input         auto_in_e_valid,
  input         auto_in_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [2:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [2:0]  auto_out_c_bits_size,
  output [6:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [2:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output        auto_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_bits_sink; // @[Nodes.scala 24:25]
  wire  a_repeater_clock; // @[HintHandler.scala 53:30]
  wire  a_repeater_reset; // @[HintHandler.scala 53:30]
  wire  a_repeater_io_repeat; // @[HintHandler.scala 53:30]
  wire  a_repeater_io_full; // @[HintHandler.scala 53:30]
  wire  a_repeater_io_enq_ready; // @[HintHandler.scala 53:30]
  wire  a_repeater_io_enq_valid; // @[HintHandler.scala 53:30]
  wire [2:0] a_repeater_io_enq_bits_size; // @[HintHandler.scala 53:30]
  wire [5:0] a_repeater_io_enq_bits_source; // @[HintHandler.scala 53:30]
  wire [31:0] a_repeater_io_enq_bits_address; // @[HintHandler.scala 53:30]
  wire  a_repeater_io_deq_ready; // @[HintHandler.scala 53:30]
  wire  a_repeater_io_deq_valid; // @[HintHandler.scala 53:30]
  wire [2:0] a_repeater_io_deq_bits_size; // @[HintHandler.scala 53:30]
  wire [5:0] a_repeater_io_deq_bits_source; // @[HintHandler.scala 53:30]
  wire [31:0] a_repeater_io_deq_bits_address; // @[HintHandler.scala 53:30]
  wire  isHint = auto_in_a_bits_opcode == 3'h5; // @[HintHandler.scala 35:37]
  wire [31:0] _helpPP_T = auto_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _helpPP_T_1 = {1'b0,$signed(_helpPP_T)}; // @[Parameters.scala 137:49]
  wire [32:0] _helpPP_T_3 = $signed(_helpPP_T_1) & 33'shf0000000; // @[Parameters.scala 137:52]
  wire  _helpPP_T_4 = $signed(_helpPP_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _helpPP_T_5 = auto_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _helpPP_T_6 = {1'b0,$signed(_helpPP_T_5)}; // @[Parameters.scala 137:49]
  wire [32:0] _helpPP_T_8 = $signed(_helpPP_T_6) & 33'she0000000; // @[Parameters.scala 137:52]
  wire  _helpPP_T_9 = $signed(_helpPP_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _helpPP_T_10 = auto_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _helpPP_T_11 = {1'b0,$signed(_helpPP_T_10)}; // @[Parameters.scala 137:49]
  wire [32:0] _helpPP_T_13 = $signed(_helpPP_T_11) & 33'shc0000000; // @[Parameters.scala 137:52]
  wire  _helpPP_T_14 = $signed(_helpPP_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _helpPP_T_15 = auto_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _helpPP_T_16 = {1'b0,$signed(_helpPP_T_15)}; // @[Parameters.scala 137:49]
  wire [32:0] _helpPP_T_18 = $signed(_helpPP_T_16) & 33'shc0000000; // @[Parameters.scala 137:52]
  wire  _helpPP_T_19 = $signed(_helpPP_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _helpPP_T_20 = auto_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _helpPP_T_21 = {1'b0,$signed(_helpPP_T_20)}; // @[Parameters.scala 137:49]
  wire [32:0] _helpPP_T_23 = $signed(_helpPP_T_21) & 33'she0000000; // @[Parameters.scala 137:52]
  wire  _helpPP_T_24 = $signed(_helpPP_T_23) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _helpPP_T_28 = _helpPP_T_4 | _helpPP_T_9 | _helpPP_T_14 | _helpPP_T_19 | _helpPP_T_24; // @[Parameters.scala 615:89]
  wire  helpPP = isHint & _helpPP_T_28; // @[HintHandler.scala 40:27]
  wire  a_valid = a_repeater_io_deq_valid; // @[HintHandler.scala 54:23 HintHandler.scala 75:19]
  wire  _a_repeater_io_repeat_T = auto_out_a_ready & a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] a_bits_size = a_repeater_io_deq_bits_size; // @[HintHandler.scala 54:23 HintHandler.scala 63:26]
  wire [12:0] _a_repeater_io_repeat_beats1_decode_T_1 = 13'h3f << a_bits_size; // @[package.scala 234:77]
  wire [5:0] _a_repeater_io_repeat_beats1_decode_T_3 = ~_a_repeater_io_repeat_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] a_repeater_io_repeat_beats1_decode = _a_repeater_io_repeat_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  mapPP = a_repeater_io_full | helpPP; // @[HintHandler.scala 78:35]
  wire [2:0] bundleOut_0_a_bits_opcode = mapPP ? 3'h1 : auto_in_a_bits_opcode; // @[HintHandler.scala 83:31]
  wire  a_repeater_io_repeat_beats1_opdata = ~bundleOut_0_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] a_repeater_io_repeat_beats1 = a_repeater_io_repeat_beats1_opdata ? a_repeater_io_repeat_beats1_decode : 3'h0
    ; // @[Edges.scala 220:14]
  reg [2:0] a_repeater_io_repeat_counter; // @[Edges.scala 228:27]
  wire [2:0] a_repeater_io_repeat_counter1 = a_repeater_io_repeat_counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_repeater_io_repeat_first = a_repeater_io_repeat_counter == 3'h0; // @[Edges.scala 230:25]
  wire  a_repeater_io_repeat_last = a_repeater_io_repeat_counter == 3'h1 | a_repeater_io_repeat_beats1 == 3'h0; // @[Edges.scala 231:37]
  wire [5:0] a_bits_source = a_repeater_io_deq_bits_source; // @[HintHandler.scala 54:23 HintHandler.scala 64:26]
  wire [6:0] _bundleOut_0_a_bits_source_T = {a_bits_source, 1'h0}; // @[HintHandler.scala 86:42]
  wire [6:0] _GEN_1 = {{6'd0}, mapPP}; // @[HintHandler.scala 86:47]
  wire  transform = auto_out_d_bits_source[0]; // @[HintHandler.scala 94:40]
  TLMonitor_14 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_c_ready(monitor_io_in_c_ready),
    .io_in_c_valid(monitor_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_io_in_c_bits_address),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),
    .io_in_e_ready(monitor_io_in_e_ready),
    .io_in_e_valid(monitor_io_in_e_valid),
    .io_in_e_bits_sink(monitor_io_in_e_bits_sink)
  );
  Repeater_1 a_repeater ( // @[HintHandler.scala 53:30]
    .clock(a_repeater_clock),
    .reset(a_repeater_reset),
    .io_repeat(a_repeater_io_repeat),
    .io_full(a_repeater_io_full),
    .io_enq_ready(a_repeater_io_enq_ready),
    .io_enq_valid(a_repeater_io_enq_valid),
    .io_enq_bits_size(a_repeater_io_enq_bits_size),
    .io_enq_bits_source(a_repeater_io_enq_bits_source),
    .io_enq_bits_address(a_repeater_io_enq_bits_address),
    .io_deq_ready(a_repeater_io_deq_ready),
    .io_deq_valid(a_repeater_io_deq_valid),
    .io_deq_bits_size(a_repeater_io_deq_bits_size),
    .io_deq_bits_source(a_repeater_io_deq_bits_source),
    .io_deq_bits_address(a_repeater_io_deq_bits_address)
  );
  assign auto_in_a_ready = a_repeater_io_enq_ready; // @[Nodes.scala 1210:84 BundleMap.scala 247:19]
  assign auto_in_c_ready = auto_out_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[HintHandler.scala 104:33]
  assign auto_in_d_bits_opcode = transform ? 3'h2 : auto_out_d_bits_opcode; // @[HintHandler.scala 103:30]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source[6:1]; // @[HintHandler.scala 102:45]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_e_ready = auto_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = a_repeater_io_deq_valid; // @[HintHandler.scala 54:23 HintHandler.scala 75:19]
  assign auto_out_a_bits_opcode = mapPP ? 3'h1 : auto_in_a_bits_opcode; // @[HintHandler.scala 83:31]
  assign auto_out_a_bits_param = mapPP ? 3'h0 : auto_in_a_bits_param; // @[HintHandler.scala 84:31]
  assign auto_out_a_bits_size = a_repeater_io_deq_bits_size; // @[HintHandler.scala 54:23 HintHandler.scala 63:26]
  assign auto_out_a_bits_source = _bundleOut_0_a_bits_source_T | _GEN_1; // @[HintHandler.scala 86:47]
  assign auto_out_a_bits_address = a_repeater_io_deq_bits_address; // @[HintHandler.scala 54:23 HintHandler.scala 65:26]
  assign auto_out_a_bits_mask = mapPP ? 8'h0 : auto_in_a_bits_mask; // @[HintHandler.scala 85:31]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_source = {auto_in_c_bits_source, 1'h0}; // @[HintHandler.scala 109:47]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[HintHandler.scala 105:33]
  assign auto_out_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = a_repeater_io_enq_ready; // @[Nodes.scala 1210:84 BundleMap.scala 247:19]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_ready = auto_out_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = auto_out_d_valid; // @[HintHandler.scala 104:33]
  assign monitor_io_in_d_bits_opcode = transform ? 3'h2 : auto_out_d_bits_opcode; // @[HintHandler.scala 103:30]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source[6:1]; // @[HintHandler.scala 102:45]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_e_ready = auto_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_repeater_clock = clock;
  assign a_repeater_reset = reset;
  assign a_repeater_io_repeat = mapPP & ~a_repeater_io_repeat_last; // @[HintHandler.scala 56:37]
  assign a_repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_repeater_io_repeat_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_repeater_io_repeat_T) begin // @[Edges.scala 234:17]
      if (a_repeater_io_repeat_first) begin // @[Edges.scala 235:21]
        if (a_repeater_io_repeat_beats1_opdata) begin // @[Edges.scala 220:14]
          a_repeater_io_repeat_counter <= a_repeater_io_repeat_beats1_decode;
        end else begin
          a_repeater_io_repeat_counter <= 3'h0;
        end
      end else begin
        a_repeater_io_repeat_counter <= a_repeater_io_repeat_counter1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_repeater_io_repeat_counter = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_15(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [5:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [3:0]  io_in_a_bits_mask,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [2:0]  io_in_c_bits_size,
  input  [5:0]  io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [5:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input         io_in_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [255:0] _RAND_19;
  reg [255:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [255:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_86 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_lo_lo = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_lo_hi = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_hi_lo = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_hi_hi = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire [31:0] _T_180 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_181 = {1'b0,$signed(_T_180)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_183 = $signed(_T_181) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_184 = $signed(_T_183) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_185 = io_in_a_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_186 = {1'b0,$signed(_T_185)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_188 = $signed(_T_186) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_189 = $signed(_T_188) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_190 = io_in_a_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_191 = {1'b0,$signed(_T_190)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_193 = $signed(_T_191) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_194 = $signed(_T_193) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_195 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_196 = {1'b0,$signed(_T_195)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_198 = $signed(_T_196) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _T_199 = $signed(_T_198) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _T_200 = io_in_a_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _T_201 = {1'b0,$signed(_T_200)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_203 = $signed(_T_201) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _T_204 = $signed(_T_203) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_211 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [31:0] _T_214 = io_in_a_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _T_215 = {1'b0,$signed(_T_214)}; // @[Parameters.scala 137:49]
  wire [32:0] _T_217 = $signed(_T_215) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _T_218 = $signed(_T_217) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _T_219 = _T_211 & _T_218; // @[Parameters.scala 670:56]
  wire  _T_222 = source_ok & _T_219; // @[Monitor.scala 82:72]
  wire  _T_277 = _source_ok_T_1 & _T_211; // @[Mux.scala 27:72]
  wire  _T_330 = _T_218 | _T_184 | _T_189 | _T_194 | _T_199 | _T_204; // @[Parameters.scala 671:42]
  wire  _T_333 = _T_277 & _T_330; // @[Monitor.scala 83:78]
  wire  _T_347 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [3:0] _T_351 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_352 = _T_351 == 4'h0; // @[Monitor.scala 88:31]
  wire  _T_360 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_593 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_606 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_709 = _T_211 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_720 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_724 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_732 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_834 = source_ok & _T_709; // @[Monitor.scala 115:71]
  wire  _T_852 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [3:0] _T_968 = ~mask; // @[Monitor.scala 127:33]
  wire [3:0] _T_969 = io_in_a_bits_mask & _T_968; // @[Monitor.scala 127:31]
  wire  _T_970 = _T_969 == 4'h0; // @[Monitor.scala 127:40]
  wire  _T_974 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_1036 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 92:42]
  wire  _T_1074 = _T_1036 & _T_330; // @[Parameters.scala 670:56]
  wire  _T_1076 = source_ok & _T_1074; // @[Monitor.scala 131:74]
  wire  _T_1086 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_1094 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_1206 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_1214 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1326 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1338 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1342 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1346 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27]
  wire  _T_1350 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_1354 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1358 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1362 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1373 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_1377 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_1390 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1410 = _T_1358 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1419 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1436 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1454 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _source_ok_T_109 = io_in_c_bits_source[5:3] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_115 = io_in_c_bits_source[5:3] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_121 = io_in_c_bits_source[5:3] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_127 = io_in_c_bits_source[5:3] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_133 = io_in_c_bits_source[5:3] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_139 = io_in_c_bits_source[5:3] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_145 = io_in_c_bits_source[5:3] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_151 = io_in_c_bits_source[5:3] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_2 = _source_ok_T_109 | _source_ok_T_115 | _source_ok_T_121 | _source_ok_T_127 | _source_ok_T_133 |
    _source_ok_T_139 | _source_ok_T_145 | _source_ok_T_151; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_7 = 13'h3f << io_in_c_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask_2 = ~_is_aligned_mask_T_7[5:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_87 = {{26'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T_2 = io_in_c_bits_address & _GEN_87; // @[Edges.scala 20:16]
  wire  is_aligned_2 = _is_aligned_T_2 == 32'h0; // @[Edges.scala 20:24]
  wire [31:0] _address_ok_T_34 = io_in_c_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_35 = {1'b0,$signed(_address_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_37 = $signed(_address_ok_T_35) & -33'sh10000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_38 = $signed(_address_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_39 = io_in_c_bits_address ^ 32'h20000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_40 = {1'b0,$signed(_address_ok_T_39)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_42 = $signed(_address_ok_T_40) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_43 = $signed(_address_ok_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_44 = io_in_c_bits_address ^ 32'h40000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_45 = {1'b0,$signed(_address_ok_T_44)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_47 = $signed(_address_ok_T_45) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_48 = $signed(_address_ok_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_49 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_50 = {1'b0,$signed(_address_ok_T_49)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_52 = $signed(_address_ok_T_50) & -33'sh40000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_53 = $signed(_address_ok_T_52) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_54 = io_in_c_bits_address ^ 32'hc0000000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_55 = {1'b0,$signed(_address_ok_T_54)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_57 = $signed(_address_ok_T_55) & -33'sh20000000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_58 = $signed(_address_ok_T_57) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _address_ok_T_62 = _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 | _address_ok_T_58; // @[Parameters.scala 598:92]
  wire [31:0] _address_ok_T_63 = io_in_c_bits_address ^ 32'h1000; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_64 = {1'b0,$signed(_address_ok_T_63)}; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_66 = $signed(_address_ok_T_64) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_67 = $signed(_address_ok_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  wire  address_ok_1 = _address_ok_T_62 | _address_ok_T_67; // @[Parameters.scala 622:64]
  wire  _T_2224 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  wire  _T_2231 = io_in_c_bits_size >= 3'h2; // @[Monitor.scala 245:30]
  wire  _T_2238 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  wire  _T_2246 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  wire  _T_2264 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  wire  _T_2357 = io_in_c_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_2365 = _T_2357 & _address_ok_T_67; // @[Parameters.scala 670:56]
  wire  _T_2368 = source_ok_2 & _T_2365; // @[Monitor.scala 260:78]
  wire  _T_2423 = _source_ok_T_109 & _T_2357; // @[Mux.scala 27:72]
  wire  _T_2476 = _address_ok_T_67 | _address_ok_T_38 | _address_ok_T_43 | _address_ok_T_48 | _address_ok_T_53 |
    _address_ok_T_58; // @[Parameters.scala 671:42]
  wire  _T_2479 = _T_2423 & _T_2476; // @[Monitor.scala 261:78]
  wire  _T_2501 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  wire  _T_2734 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  wire  _T_2744 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  wire  _T_2752 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  wire  _T_2766 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  wire  sink_ok_1 = io_in_e_bits_sink < 1'h1; // @[Monitor.scala 364:31]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [5:0] source; // @[Monitor.scala 387:22]
  reg [31:0] address; // @[Monitor.scala 388:22]
  wire  _T_2788 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_2789 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_2793 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_2797 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_2801 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_2805 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [5:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_2812 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_2813 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_2817 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_2821 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_2825 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_2833 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  wire  _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  wire [3:0] c_first_beats1_decode = is_aligned_mask_2[5:2]; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  reg [3:0] c_first_counter; // @[Edges.scala 228:27]
  wire [3:0] c_first_counter1 = c_first_counter - 4'h1; // @[Edges.scala 229:28]
  wire  c_first = c_first_counter == 4'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [2:0] size_3; // @[Monitor.scala 514:22]
  reg [5:0] source_3; // @[Monitor.scala 515:22]
  reg [31:0] address_2; // @[Monitor.scala 516:22]
  wire  _T_2864 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  wire  _T_2865 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  wire  _T_2869 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  wire  _T_2873 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  wire  _T_2877 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  wire  _T_2881 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  reg [63:0] inflight; // @[Monitor.scala 611:27]
  reg [255:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [255:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  wire [7:0] _GEN_88 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [8:0] _a_opcode_lookup_T = {{1'd0}, _GEN_88}; // @[Monitor.scala 634:69]
  wire [255:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [255:0] _GEN_89 = {{240'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [255:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_89; // @[Monitor.scala 634:97]
  wire [255:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[255:1]}; // @[Monitor.scala 634:152]
  wire [255:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [255:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 638:91]
  wire [255:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[255:1]}; // @[Monitor.scala 638:144]
  wire  _T_2887 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [63:0] _a_set_wo_ready_T = 64'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 64'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_2890 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [7:0] _GEN_94 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [8:0] _a_opcodes_set_T = {{1'd0}, _GEN_94}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [514:0] _GEN_95 = {{511'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [514:0] _a_opcodes_set_T_1 = _GEN_95 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [514:0] _GEN_97 = {{511'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [514:0] _a_sizes_set_T_1 = _GEN_97 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [63:0] _T_2892 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_2894 = ~_T_2892[0]; // @[Monitor.scala 658:17]
  wire [63:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 64'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [514:0] _GEN_31 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 515'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [514:0] _GEN_32 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 515'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_2898 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_2900 = ~_T_1342; // @[Monitor.scala 671:74]
  wire  _T_2901 = io_in_d_valid & d_first_1 & ~_T_1342; // @[Monitor.scala 671:71]
  wire [63:0] _d_clr_wo_ready_T = 64'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [526:0] _GEN_99 = {{511'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [526:0] _d_opcodes_clr_T_5 = _GEN_99 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [63:0] d_clr = _d_first_T & d_first_1 & _T_2900 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [526:0] _GEN_35 = _d_first_T & d_first_1 & _T_2900 ? _d_opcodes_clr_T_5 : 527'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_2887 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [63:0] _T_2911 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_2913 = _T_2911[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_2918 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_2919 = io_in_d_bits_opcode == _GEN_44 | _T_2918; // @[Monitor.scala 685:77]
  wire  _T_2923 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_2930 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_2931 = io_in_d_bits_opcode == _GEN_60 | _T_2930; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_102 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_2935 = _GEN_102 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_2945 = _T_2898 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_2900; // @[Monitor.scala 694:116]
  wire  _T_2946 = ~io_in_d_ready; // @[Monitor.scala 695:15]
  wire  _T_2947 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_2954 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [63:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [63:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [63:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [255:0] a_opcodes_set = _GEN_31[255:0];
  wire [255:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [255:0] d_opcodes_clr = _GEN_35[255:0];
  wire [255:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [255:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [255:0] a_sizes_set = _GEN_32[255:0];
  wire [255:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [255:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_2963 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [63:0] inflight_1; // @[Monitor.scala 723:35]
  reg [255:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [3:0] c_first_counter_1; // @[Edges.scala 228:27]
  wire [3:0] c_first_counter1_1 = c_first_counter_1 - 4'h1; // @[Edges.scala 229:28]
  wire  c_first_1 = c_first_counter_1 == 4'h0; // @[Edges.scala 230:25]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25]
  wire [255:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [255:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 747:93]
  wire [255:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[255:1]}; // @[Monitor.scala 747:146]
  wire  _T_2973 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  _T_2974 = io_in_c_valid & c_first_1 & _T_2973; // @[Monitor.scala 756:37]
  wire [63:0] _c_set_wo_ready_T = 64'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  wire [63:0] c_set_wo_ready = io_in_c_valid & c_first_1 & _T_2973 ? _c_set_wo_ready_T : 64'h0; // @[Monitor.scala 756:71 Monitor.scala 757:22]
  wire  _T_2980 = _c_first_T & c_first_1 & _T_2973; // @[Monitor.scala 760:38]
  wire [3:0] _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  wire [3:0] _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 4'h1; // @[Monitor.scala 763:59]
  wire [7:0] _GEN_109 = {io_in_c_bits_source, 2'h0}; // @[Monitor.scala 764:79]
  wire [8:0] _c_opcodes_set_T = {{1'd0}, _GEN_109}; // @[Monitor.scala 764:79]
  wire [3:0] c_sizes_set_interm = _c_first_T & c_first_1 & _T_2973 ? _c_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 760:72 Monitor.scala 763:28]
  wire [514:0] _GEN_112 = {{511'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  wire [514:0] _c_sizes_set_T_1 = _GEN_112 << _c_opcodes_set_T; // @[Monitor.scala 765:52]
  wire [63:0] _T_2981 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  wire  _T_2983 = ~_T_2981[0]; // @[Monitor.scala 766:17]
  wire [63:0] c_set = _c_first_T & c_first_1 & _T_2973 ? _c_set_wo_ready_T : 64'h0; // @[Monitor.scala 760:72 Monitor.scala 761:28]
  wire [514:0] _GEN_77 = _c_first_T & c_first_1 & _T_2973 ? _c_sizes_set_T_1 : 515'h0; // @[Monitor.scala 760:72 Monitor.scala 765:28]
  wire  _T_2987 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  wire  _T_2989 = io_in_d_valid & d_first_2 & _T_1342; // @[Monitor.scala 779:71]
  wire [63:0] d_clr_wo_ready_1 = io_in_d_valid & d_first_2 & _T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 779:89 Monitor.scala 780:22]
  wire [63:0] d_clr_1 = _d_first_T & d_first_2 & _T_1342 ? _d_clr_wo_ready_T : 64'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [526:0] _GEN_80 = _d_first_T & d_first_2 & _T_1342 ? _d_opcodes_clr_T_5 : 527'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire  _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1 = _T_2974 & io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:88]
  wire [63:0] _T_2997 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire  _T_2999 = _T_2997[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  wire  _T_3003 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_3007 = _GEN_102 == c_size_lookup; // @[Monitor.scala 795:36]
  wire  _T_3016 = _T_2987 & c_first_1 & io_in_c_valid & _same_cycle_resp_T_8 & _T_1342; // @[Monitor.scala 799:116]
  wire  _T_3018 = _T_2946 | io_in_c_ready; // @[Monitor.scala 800:32]
  wire  _T_3022 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  wire  _T_3023 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  wire [63:0] _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  wire [63:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [63:0] _inflight_T_5 = _inflight_T_3 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [255:0] d_opcodes_clr_1 = _GEN_80[255:0];
  wire [255:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [255:0] c_sizes_set = _GEN_77[255:0];
  wire [255:0] _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  wire [255:0] _inflight_sizes_T_5 = _inflight_sizes_T_3 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_3032 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [3:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [3:0] d_first_counter1_3 = d_first_counter_3 - 4'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 4'h0; // @[Edges.scala 230:25]
  wire  _T_3044 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_3045 = _d_first_T & d_first_3 & _T_3044; // @[Monitor.scala 829:38]
  wire  _T_3048 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = _d_first_T & d_first_3 & _T_3044 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  _T_3052 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _e_clr_T = 2'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  wire  d_set = _GEN_84[0];
  wire  _T_3056 = (d_set | inflight_2) >> io_in_e_bits_sink; // @[Monitor.scala 837:35]
  wire [1:0] _GEN_85 = _T_3052 ? _e_clr_T : 2'h0; // @[Monitor.scala 835:73 Monitor.scala 836:13]
  wire  e_clr = _GEN_85[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter <= 4'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 4'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      opcode_3 <= io_in_c_bits_opcode; // @[Monitor.scala 525:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      param_3 <= io_in_c_bits_param; // @[Monitor.scala 526:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      size_3 <= io_in_c_bits_size; // @[Monitor.scala 527:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      source_3 <= io_in_c_bits_source; // @[Monitor.scala 528:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      address_2 <= io_in_c_bits_address; // @[Monitor.scala 529:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 64'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 256'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 256'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 64'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 256'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter_1 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first_1) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 4'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_c_first_T | _d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= (inflight_2 | d_set) & ~e_clr; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 4'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 4'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_222 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_333 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_347 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_593 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_360 & ~(_T_352 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_709 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_606 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_732 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_720 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_852 & ~(_T_970 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_1086 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_974 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1076 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_1206 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1094 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_834 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_834 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1326 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_1326 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_1214 & ~(_T_724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1338 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1338 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1358 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1342 & ~(_T_1358 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1373 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1373 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1377 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1377 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1362 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1346 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1346 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1373 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1373 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1377 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1377 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1390 & ~(_T_1410 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1419 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1436 & ~(_T_1410 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1350 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1350 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1354 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1454 & ~(_T_1354 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2224 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2246 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2368 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2368 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2479 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2479 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid report param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2264 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2368 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2368 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2479 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2479 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2238 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2501 & ~(_T_2238 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2734 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2752 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(address_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(address_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(_T_2744 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2766 & ~(_T_2744 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channels carries invalid sink ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & ~(sink_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2789 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2789 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2793 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2793 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2797 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2797 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2801 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2801 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2788 & ~(_T_2805 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2788 & ~(_T_2805 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2813 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2813 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2817 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2817 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2821 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2821 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2825 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2825 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2812 & ~(_T_2833 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2812 & ~(_T_2833 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2865 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2865 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2869 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2869 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2873 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2873 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2877 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2877 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2864 & ~(_T_2881 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2864 & ~(_T_2881 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2890 & ~(_T_2894 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2890 & ~(_T_2894 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~(_T_2913 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~(_T_2913 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2919 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2919 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2923 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & same_cycle_resp & ~(_T_2923 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2931 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2931 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2935 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901 & ~same_cycle_resp & ~(_T_2935 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2945 & ~(_T_2947 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2945 & ~(_T_2947 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2954 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2954 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2963 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2963 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2980 & ~(_T_2983 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel re-used a source ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2980 & ~(_T_2983 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & ~(_T_2999 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & ~(_T_2999 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & same_cycle_resp_1 & ~(_T_3003 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & same_cycle_resp_1 & ~(_T_3003 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2989 & ~same_cycle_resp_1 & ~(_T_3007 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2989 & ~same_cycle_resp_1 & ~(_T_3007 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3016 & ~(_T_3018 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3016 & ~(_T_3018 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3022 & ~(_T_3023 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3022 & ~(_T_3023 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_3032 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_3032 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3045 & ~(_T_3048 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3045 & ~(_T_3048 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3052 & ~(_T_3056 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:153:118)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3052 & ~(_T_3056 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  c_first_counter = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  opcode_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  param_3 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  size_3 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  source_3 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  address_2 = _RAND_17[31:0];
  _RAND_18 = {2{`RANDOM}};
  inflight = _RAND_18[63:0];
  _RAND_19 = {8{`RANDOM}};
  inflight_opcodes = _RAND_19[255:0];
  _RAND_20 = {8{`RANDOM}};
  inflight_sizes = _RAND_20[255:0];
  _RAND_21 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  watchdog = _RAND_23[31:0];
  _RAND_24 = {2{`RANDOM}};
  inflight_1 = _RAND_24[63:0];
  _RAND_25 = {8{`RANDOM}};
  inflight_sizes_1 = _RAND_25[255:0];
  _RAND_26 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  watchdog_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inflight_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_30[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_2(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [5:0]  io_enq_bits_source,
  input         io_enq_bits_denied,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [5:0]  io_deq_bits_source,
  output        io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [1:0] saved_param; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [5:0] saved_source; // @[Repeater.scala 20:18]
  reg  saved_denied; // @[Repeater.scala 20:18]
  reg [63:0] saved_data; // @[Repeater.scala 20:18]
  reg  saved_corrupt; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 28:38 Repeater.scala 28:45 Repeater.scala 19:21]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_denied = full ? saved_denied : io_enq_bits_denied; // @[Repeater.scala 25:21]
  assign io_deq_bits_data = full ? saved_data : io_enq_bits_data; // @[Repeater.scala 25:21]
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; // @[Repeater.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin // @[Repeater.scala 29:38]
      full <= 1'h0; // @[Repeater.scala 29:45]
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_param <= io_enq_bits_param; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_denied <= io_enq_bits_denied; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_data <= io_enq_bits_data; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_corrupt <= io_enq_bits_corrupt; // @[Repeater.scala 28:62]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  saved_denied = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  saved_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  saved_corrupt = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLWidthWidget_1(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [5:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [3:0]  auto_in_a_bits_mask,
  input  [31:0] auto_in_a_bits_data,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [2:0]  auto_in_c_bits_size,
  input  [5:0]  auto_in_c_bits_source,
  input  [31:0] auto_in_c_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [5:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [31:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  output        auto_in_e_ready,
  input         auto_in_e_valid,
  input         auto_in_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [2:0]  auto_out_a_bits_size,
  output [5:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [2:0]  auto_out_c_bits_size,
  output [5:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [2:0]  auto_out_d_bits_size,
  input  [5:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output        auto_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [5:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_bits_sink; // @[Nodes.scala 24:25]
  wire  repeated_repeater_clock; // @[Repeater.scala 35:26]
  wire  repeated_repeater_reset; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_repeat; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_opcode; // @[Repeater.scala 35:26]
  wire [1:0] repeated_repeater_io_enq_bits_param; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_size; // @[Repeater.scala 35:26]
  wire [5:0] repeated_repeater_io_enq_bits_source; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_bits_denied; // @[Repeater.scala 35:26]
  wire [63:0] repeated_repeater_io_enq_bits_data; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_bits_corrupt; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_opcode; // @[Repeater.scala 35:26]
  wire [1:0] repeated_repeater_io_deq_bits_param; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_size; // @[Repeater.scala 35:26]
  wire [5:0] repeated_repeater_io_deq_bits_source; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_bits_denied; // @[Repeater.scala 35:26]
  wire [63:0] repeated_repeater_io_deq_bits_data; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_bits_corrupt; // @[Repeater.scala 35:26]
  wire  hasData = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [9:0] _limit_T_1 = 10'h7 << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [2:0] _limit_T_3 = ~_limit_T_1[2:0]; // @[package.scala 234:46]
  wire  limit = _limit_T_3[2]; // @[WidthWidget.scala 32:47]
  reg  count; // @[WidthWidget.scala 34:27]
  wire  last = count == limit | ~hasData; // @[WidthWidget.scala 36:36]
  wire  enable_0 = ~(|(count & limit)); // @[WidthWidget.scala 37:47]
  wire  _bundleIn_0_a_ready_T = ~last; // @[WidthWidget.scala 70:32]
  wire  bundleIn_0_a_ready = auto_out_a_ready | ~last; // @[WidthWidget.scala 70:29]
  wire  _T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37]
  reg  bundleOut_0_a_bits_data_rdata_written_once; // @[WidthWidget.scala 56:41]
  wire  bundleOut_0_a_bits_data_masked_enable_0 = enable_0 | ~bundleOut_0_a_bits_data_rdata_written_once; // @[WidthWidget.scala 57:42]
  reg [31:0] bundleOut_0_a_bits_data_rdata_0; // @[WidthWidget.scala 60:24]
  wire [31:0] bundleOut_0_a_bits_data_lo = bundleOut_0_a_bits_data_masked_enable_0 ? auto_in_a_bits_data :
    bundleOut_0_a_bits_data_rdata_0; // @[WidthWidget.scala 62:88]
  wire  _GEN_4 = _T & _bundleIn_0_a_ready_T | bundleOut_0_a_bits_data_rdata_written_once; // @[WidthWidget.scala 63:35 WidthWidget.scala 64:30 WidthWidget.scala 56:41]
  wire [1:0] bundleOut_0_a_bits_mask_sizeOH_shiftAmount = auto_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _bundleOut_0_a_bits_mask_sizeOH_T_1 = 4'h1 << bundleOut_0_a_bits_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] bundleOut_0_a_bits_mask_sizeOH = _bundleOut_0_a_bits_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _bundleOut_0_a_bits_mask_T = auto_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  bundleOut_0_a_bits_mask_size = bundleOut_0_a_bits_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  bundleOut_0_a_bits_mask_bit = auto_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  bundleOut_0_a_bits_mask_nbit = ~bundleOut_0_a_bits_mask_bit; // @[Misc.scala 210:20]
  wire  bundleOut_0_a_bits_mask_acc = _bundleOut_0_a_bits_mask_T | bundleOut_0_a_bits_mask_size &
    bundleOut_0_a_bits_mask_nbit; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_acc_1 = _bundleOut_0_a_bits_mask_T | bundleOut_0_a_bits_mask_size &
    bundleOut_0_a_bits_mask_bit; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_size_1 = bundleOut_0_a_bits_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  bundleOut_0_a_bits_mask_bit_1 = auto_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  bundleOut_0_a_bits_mask_nbit_1 = ~bundleOut_0_a_bits_mask_bit_1; // @[Misc.scala 210:20]
  wire  bundleOut_0_a_bits_mask_eq_2 = bundleOut_0_a_bits_mask_nbit & bundleOut_0_a_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_acc_2 = bundleOut_0_a_bits_mask_acc | bundleOut_0_a_bits_mask_size_1 &
    bundleOut_0_a_bits_mask_eq_2; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_3 = bundleOut_0_a_bits_mask_nbit & bundleOut_0_a_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_acc_3 = bundleOut_0_a_bits_mask_acc | bundleOut_0_a_bits_mask_size_1 &
    bundleOut_0_a_bits_mask_eq_3; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_4 = bundleOut_0_a_bits_mask_bit & bundleOut_0_a_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_acc_4 = bundleOut_0_a_bits_mask_acc_1 | bundleOut_0_a_bits_mask_size_1 &
    bundleOut_0_a_bits_mask_eq_4; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_5 = bundleOut_0_a_bits_mask_bit & bundleOut_0_a_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_acc_5 = bundleOut_0_a_bits_mask_acc_1 | bundleOut_0_a_bits_mask_size_1 &
    bundleOut_0_a_bits_mask_eq_5; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_size_2 = bundleOut_0_a_bits_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  bundleOut_0_a_bits_mask_bit_2 = auto_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  bundleOut_0_a_bits_mask_nbit_2 = ~bundleOut_0_a_bits_mask_bit_2; // @[Misc.scala 210:20]
  wire  bundleOut_0_a_bits_mask_eq_6 = bundleOut_0_a_bits_mask_eq_2 & bundleOut_0_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_lo_lo_lo = bundleOut_0_a_bits_mask_acc_2 | bundleOut_0_a_bits_mask_size_2 &
    bundleOut_0_a_bits_mask_eq_6; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_7 = bundleOut_0_a_bits_mask_eq_2 & bundleOut_0_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_lo_lo_hi = bundleOut_0_a_bits_mask_acc_2 | bundleOut_0_a_bits_mask_size_2 &
    bundleOut_0_a_bits_mask_eq_7; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_8 = bundleOut_0_a_bits_mask_eq_3 & bundleOut_0_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_lo_hi_lo = bundleOut_0_a_bits_mask_acc_3 | bundleOut_0_a_bits_mask_size_2 &
    bundleOut_0_a_bits_mask_eq_8; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_9 = bundleOut_0_a_bits_mask_eq_3 & bundleOut_0_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_lo_hi_hi = bundleOut_0_a_bits_mask_acc_3 | bundleOut_0_a_bits_mask_size_2 &
    bundleOut_0_a_bits_mask_eq_9; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_10 = bundleOut_0_a_bits_mask_eq_4 & bundleOut_0_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_hi_lo_lo = bundleOut_0_a_bits_mask_acc_4 | bundleOut_0_a_bits_mask_size_2 &
    bundleOut_0_a_bits_mask_eq_10; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_11 = bundleOut_0_a_bits_mask_eq_4 & bundleOut_0_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_hi_lo_hi = bundleOut_0_a_bits_mask_acc_4 | bundleOut_0_a_bits_mask_size_2 &
    bundleOut_0_a_bits_mask_eq_11; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_12 = bundleOut_0_a_bits_mask_eq_5 & bundleOut_0_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_hi_hi_lo = bundleOut_0_a_bits_mask_acc_5 | bundleOut_0_a_bits_mask_size_2 &
    bundleOut_0_a_bits_mask_eq_12; // @[Misc.scala 214:29]
  wire  bundleOut_0_a_bits_mask_eq_13 = bundleOut_0_a_bits_mask_eq_5 & bundleOut_0_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  bundleOut_0_a_bits_mask_hi_hi_hi = bundleOut_0_a_bits_mask_acc_5 | bundleOut_0_a_bits_mask_size_2 &
    bundleOut_0_a_bits_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] _bundleOut_0_a_bits_mask_T_1 = {bundleOut_0_a_bits_mask_hi_hi_hi,bundleOut_0_a_bits_mask_hi_hi_lo,
    bundleOut_0_a_bits_mask_hi_lo_hi,bundleOut_0_a_bits_mask_hi_lo_lo,bundleOut_0_a_bits_mask_lo_hi_hi,
    bundleOut_0_a_bits_mask_lo_hi_lo,bundleOut_0_a_bits_mask_lo_lo_hi,bundleOut_0_a_bits_mask_lo_lo_lo}; // @[Cat.scala 30:58]
  reg  bundleOut_0_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 56:41]
  wire  bundleOut_0_a_bits_mask_masked_enable_0 = enable_0 | ~bundleOut_0_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 57:42]
  reg [3:0] bundleOut_0_a_bits_mask_rdata_0; // @[WidthWidget.scala 60:24]
  wire [3:0] bundleOut_0_a_bits_mask_lo_1 = bundleOut_0_a_bits_mask_masked_enable_0 ? auto_in_a_bits_mask :
    bundleOut_0_a_bits_mask_rdata_0; // @[WidthWidget.scala 62:88]
  wire  _GEN_6 = _T & _bundleIn_0_a_ready_T | bundleOut_0_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 63:35 WidthWidget.scala 64:30 WidthWidget.scala 56:41]
  wire [7:0] _bundleOut_0_a_bits_mask_T_5 = {auto_in_a_bits_mask,bundleOut_0_a_bits_mask_lo_1}; // @[Cat.scala 30:58]
  wire [7:0] _bundleOut_0_a_bits_mask_T_7 = hasData ? _bundleOut_0_a_bits_mask_T_5 : 8'hff; // @[WidthWidget.scala 79:93]
  wire [31:0] cated_bits_data_hi = repeated_repeater_io_deq_bits_data[63:32]; // @[WidthWidget.scala 158:37]
  wire [31:0] cated_bits_data_lo = auto_out_d_bits_data[31:0]; // @[WidthWidget.scala 159:31]
  wire [63:0] cated_bits_data = {cated_bits_data_hi,cated_bits_data_lo}; // @[Cat.scala 30:58]
  wire [2:0] cated_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  repeat_hasData = cated_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] cated_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire [9:0] _repeat_limit_T_1 = 10'h7 << cated_bits_size; // @[package.scala 234:77]
  wire [2:0] _repeat_limit_T_3 = ~_repeat_limit_T_1[2:0]; // @[package.scala 234:46]
  wire  repeat_limit = _repeat_limit_T_3[2]; // @[WidthWidget.scala 97:47]
  reg  repeat_count; // @[WidthWidget.scala 99:26]
  wire  repeat_first = ~repeat_count; // @[WidthWidget.scala 100:25]
  wire  repeat_last = repeat_count == repeat_limit | ~repeat_hasData; // @[WidthWidget.scala 101:35]
  wire  cated_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  _repeat_T = auto_in_d_ready & cated_valid; // @[Decoupled.scala 40:37]
  reg  repeat_sel_sel_sources_0; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_1; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_2; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_3; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_4; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_5; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_6; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_7; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_8; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_9; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_10; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_11; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_12; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_13; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_14; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_15; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_16; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_17; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_18; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_19; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_20; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_21; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_22; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_23; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_24; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_25; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_26; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_27; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_28; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_29; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_30; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_31; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_32; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_33; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_34; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_35; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_36; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_37; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_38; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_39; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_40; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_41; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_42; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_43; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_44; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_45; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_46; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_47; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_48; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_49; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_50; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_51; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_52; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_53; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_54; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_55; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_56; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_57; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_58; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_59; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_60; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_61; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_62; // @[WidthWidget.scala 180:27]
  reg  repeat_sel_sel_sources_63; // @[WidthWidget.scala 180:27]
  wire [5:0] cated_bits_source = repeated_repeater_io_deq_bits_source; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  reg  repeat_sel_hold_r; // @[Reg.scala 15:16]
  wire  _GEN_139 = 6'h1 == cated_bits_source ? repeat_sel_sel_sources_1 : repeat_sel_sel_sources_0; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_140 = 6'h2 == cated_bits_source ? repeat_sel_sel_sources_2 : _GEN_139; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_141 = 6'h3 == cated_bits_source ? repeat_sel_sel_sources_3 : _GEN_140; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_142 = 6'h4 == cated_bits_source ? repeat_sel_sel_sources_4 : _GEN_141; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_143 = 6'h5 == cated_bits_source ? repeat_sel_sel_sources_5 : _GEN_142; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_144 = 6'h6 == cated_bits_source ? repeat_sel_sel_sources_6 : _GEN_143; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_145 = 6'h7 == cated_bits_source ? repeat_sel_sel_sources_7 : _GEN_144; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_146 = 6'h8 == cated_bits_source ? repeat_sel_sel_sources_8 : _GEN_145; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_147 = 6'h9 == cated_bits_source ? repeat_sel_sel_sources_9 : _GEN_146; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_148 = 6'ha == cated_bits_source ? repeat_sel_sel_sources_10 : _GEN_147; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_149 = 6'hb == cated_bits_source ? repeat_sel_sel_sources_11 : _GEN_148; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_150 = 6'hc == cated_bits_source ? repeat_sel_sel_sources_12 : _GEN_149; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_151 = 6'hd == cated_bits_source ? repeat_sel_sel_sources_13 : _GEN_150; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_152 = 6'he == cated_bits_source ? repeat_sel_sel_sources_14 : _GEN_151; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_153 = 6'hf == cated_bits_source ? repeat_sel_sel_sources_15 : _GEN_152; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_154 = 6'h10 == cated_bits_source ? repeat_sel_sel_sources_16 : _GEN_153; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_155 = 6'h11 == cated_bits_source ? repeat_sel_sel_sources_17 : _GEN_154; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_156 = 6'h12 == cated_bits_source ? repeat_sel_sel_sources_18 : _GEN_155; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_157 = 6'h13 == cated_bits_source ? repeat_sel_sel_sources_19 : _GEN_156; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_158 = 6'h14 == cated_bits_source ? repeat_sel_sel_sources_20 : _GEN_157; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_159 = 6'h15 == cated_bits_source ? repeat_sel_sel_sources_21 : _GEN_158; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_160 = 6'h16 == cated_bits_source ? repeat_sel_sel_sources_22 : _GEN_159; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_161 = 6'h17 == cated_bits_source ? repeat_sel_sel_sources_23 : _GEN_160; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_162 = 6'h18 == cated_bits_source ? repeat_sel_sel_sources_24 : _GEN_161; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_163 = 6'h19 == cated_bits_source ? repeat_sel_sel_sources_25 : _GEN_162; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_164 = 6'h1a == cated_bits_source ? repeat_sel_sel_sources_26 : _GEN_163; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_165 = 6'h1b == cated_bits_source ? repeat_sel_sel_sources_27 : _GEN_164; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_166 = 6'h1c == cated_bits_source ? repeat_sel_sel_sources_28 : _GEN_165; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_167 = 6'h1d == cated_bits_source ? repeat_sel_sel_sources_29 : _GEN_166; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_168 = 6'h1e == cated_bits_source ? repeat_sel_sel_sources_30 : _GEN_167; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_169 = 6'h1f == cated_bits_source ? repeat_sel_sel_sources_31 : _GEN_168; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_170 = 6'h20 == cated_bits_source ? repeat_sel_sel_sources_32 : _GEN_169; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_171 = 6'h21 == cated_bits_source ? repeat_sel_sel_sources_33 : _GEN_170; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_172 = 6'h22 == cated_bits_source ? repeat_sel_sel_sources_34 : _GEN_171; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_173 = 6'h23 == cated_bits_source ? repeat_sel_sel_sources_35 : _GEN_172; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_174 = 6'h24 == cated_bits_source ? repeat_sel_sel_sources_36 : _GEN_173; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_175 = 6'h25 == cated_bits_source ? repeat_sel_sel_sources_37 : _GEN_174; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_176 = 6'h26 == cated_bits_source ? repeat_sel_sel_sources_38 : _GEN_175; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_177 = 6'h27 == cated_bits_source ? repeat_sel_sel_sources_39 : _GEN_176; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_178 = 6'h28 == cated_bits_source ? repeat_sel_sel_sources_40 : _GEN_177; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_179 = 6'h29 == cated_bits_source ? repeat_sel_sel_sources_41 : _GEN_178; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_180 = 6'h2a == cated_bits_source ? repeat_sel_sel_sources_42 : _GEN_179; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_181 = 6'h2b == cated_bits_source ? repeat_sel_sel_sources_43 : _GEN_180; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_182 = 6'h2c == cated_bits_source ? repeat_sel_sel_sources_44 : _GEN_181; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_183 = 6'h2d == cated_bits_source ? repeat_sel_sel_sources_45 : _GEN_182; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_184 = 6'h2e == cated_bits_source ? repeat_sel_sel_sources_46 : _GEN_183; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_185 = 6'h2f == cated_bits_source ? repeat_sel_sel_sources_47 : _GEN_184; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_186 = 6'h30 == cated_bits_source ? repeat_sel_sel_sources_48 : _GEN_185; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_187 = 6'h31 == cated_bits_source ? repeat_sel_sel_sources_49 : _GEN_186; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_188 = 6'h32 == cated_bits_source ? repeat_sel_sel_sources_50 : _GEN_187; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_189 = 6'h33 == cated_bits_source ? repeat_sel_sel_sources_51 : _GEN_188; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_190 = 6'h34 == cated_bits_source ? repeat_sel_sel_sources_52 : _GEN_189; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_191 = 6'h35 == cated_bits_source ? repeat_sel_sel_sources_53 : _GEN_190; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_192 = 6'h36 == cated_bits_source ? repeat_sel_sel_sources_54 : _GEN_191; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_193 = 6'h37 == cated_bits_source ? repeat_sel_sel_sources_55 : _GEN_192; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_194 = 6'h38 == cated_bits_source ? repeat_sel_sel_sources_56 : _GEN_193; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_195 = 6'h39 == cated_bits_source ? repeat_sel_sel_sources_57 : _GEN_194; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_196 = 6'h3a == cated_bits_source ? repeat_sel_sel_sources_58 : _GEN_195; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_197 = 6'h3b == cated_bits_source ? repeat_sel_sel_sources_59 : _GEN_196; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_198 = 6'h3c == cated_bits_source ? repeat_sel_sel_sources_60 : _GEN_197; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_199 = 6'h3d == cated_bits_source ? repeat_sel_sel_sources_61 : _GEN_198; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_200 = 6'h3e == cated_bits_source ? repeat_sel_sel_sources_62 : _GEN_199; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_201 = 6'h3f == cated_bits_source ? repeat_sel_sel_sources_63 : _GEN_200; // @[Reg.scala 16:23 Reg.scala 16:23]
  wire  _GEN_202 = repeat_first ? _GEN_201 : repeat_sel_hold_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  wire  repeat_sel = _GEN_202 & ~repeat_limit; // @[WidthWidget.scala 116:16]
  wire  repeat_index = repeat_sel | repeat_count; // @[WidthWidget.scala 120:24]
  wire [31:0] repeat_bundleIn_0_d_bits_data_mux_0 = cated_bits_data[31:0]; // @[WidthWidget.scala 122:55]
  wire [31:0] repeat_bundleIn_0_d_bits_data_mux_1 = cated_bits_data[63:32]; // @[WidthWidget.scala 122:55]
  wire  hasData_1 = auto_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  wire [9:0] _limit_T_5 = 10'h7 << auto_in_c_bits_size; // @[package.scala 234:77]
  wire [2:0] _limit_T_7 = ~_limit_T_5[2:0]; // @[package.scala 234:46]
  wire  limit_1 = _limit_T_7[2]; // @[WidthWidget.scala 32:47]
  reg  count_1; // @[WidthWidget.scala 34:27]
  wire  last_1 = count_1 == limit_1 | ~hasData_1; // @[WidthWidget.scala 36:36]
  wire  bundleIn_0_c_ready = auto_out_c_ready | ~last_1; // @[WidthWidget.scala 70:29]
  wire  _T_1 = bundleIn_0_c_ready & auto_in_c_valid; // @[Decoupled.scala 40:37]
  TLMonitor_15 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_c_ready(monitor_io_in_c_ready),
    .io_in_c_valid(monitor_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_io_in_c_bits_address),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),
    .io_in_e_ready(monitor_io_in_e_ready),
    .io_in_e_valid(monitor_io_in_e_valid),
    .io_in_e_bits_sink(monitor_io_in_e_bits_sink)
  );
  Repeater_2 repeated_repeater ( // @[Repeater.scala 35:26]
    .clock(repeated_repeater_clock),
    .reset(repeated_repeater_reset),
    .io_repeat(repeated_repeater_io_repeat),
    .io_enq_ready(repeated_repeater_io_enq_ready),
    .io_enq_valid(repeated_repeater_io_enq_valid),
    .io_enq_bits_opcode(repeated_repeater_io_enq_bits_opcode),
    .io_enq_bits_param(repeated_repeater_io_enq_bits_param),
    .io_enq_bits_size(repeated_repeater_io_enq_bits_size),
    .io_enq_bits_source(repeated_repeater_io_enq_bits_source),
    .io_enq_bits_denied(repeated_repeater_io_enq_bits_denied),
    .io_enq_bits_data(repeated_repeater_io_enq_bits_data),
    .io_enq_bits_corrupt(repeated_repeater_io_enq_bits_corrupt),
    .io_deq_ready(repeated_repeater_io_deq_ready),
    .io_deq_valid(repeated_repeater_io_deq_valid),
    .io_deq_bits_opcode(repeated_repeater_io_deq_bits_opcode),
    .io_deq_bits_param(repeated_repeater_io_deq_bits_param),
    .io_deq_bits_size(repeated_repeater_io_deq_bits_size),
    .io_deq_bits_source(repeated_repeater_io_deq_bits_source),
    .io_deq_bits_denied(repeated_repeater_io_deq_bits_denied),
    .io_deq_bits_data(repeated_repeater_io_deq_bits_data),
    .io_deq_bits_corrupt(repeated_repeater_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = auto_out_a_ready | ~last; // @[WidthWidget.scala 70:29]
  assign auto_in_c_ready = auto_out_c_ready | ~last_1; // @[WidthWidget.scala 70:29]
  assign auto_in_d_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_in_d_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_in_d_bits_param = repeated_repeater_io_deq_bits_param; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_in_d_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_in_d_bits_source = repeated_repeater_io_deq_bits_source; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_in_d_bits_denied = repeated_repeater_io_deq_bits_denied; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_in_d_bits_data = repeat_index ? repeat_bundleIn_0_d_bits_data_mux_1 : repeat_bundleIn_0_d_bits_data_mux_0; // @[WidthWidget.scala 131:30 WidthWidget.scala 131:30]
  assign auto_in_d_bits_corrupt = repeated_repeater_io_deq_bits_corrupt; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_in_e_ready = auto_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid & last; // @[WidthWidget.scala 71:29]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = _bundleOut_0_a_bits_mask_T_1 & _bundleOut_0_a_bits_mask_T_7; // @[WidthWidget.scala 79:88]
  assign auto_out_a_bits_data = {auto_in_a_bits_data,bundleOut_0_a_bits_data_lo}; // @[Cat.scala 30:58]
  assign auto_out_c_valid = auto_in_c_valid & last_1; // @[WidthWidget.scala 71:29]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = repeated_repeater_io_enq_ready; // @[Nodes.scala 1207:84 Repeater.scala 37:21]
  assign auto_out_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = auto_out_a_ready | ~last; // @[WidthWidget.scala 70:29]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_ready = auto_out_c_ready | ~last_1; // @[WidthWidget.scala 70:29]
  assign monitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign monitor_io_in_d_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign monitor_io_in_d_bits_param = repeated_repeater_io_deq_bits_param; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign monitor_io_in_d_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign monitor_io_in_d_bits_source = repeated_repeater_io_deq_bits_source; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign monitor_io_in_d_bits_denied = repeated_repeater_io_deq_bits_denied; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign monitor_io_in_d_bits_corrupt = repeated_repeater_io_deq_bits_corrupt; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign monitor_io_in_e_ready = auto_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_e_bits_sink = auto_in_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_clock = clock;
  assign repeated_repeater_reset = reset;
  assign repeated_repeater_io_repeat = ~repeat_last; // @[WidthWidget.scala 142:7]
  assign repeated_repeater_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_io_enq_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  always @(posedge clock) begin
    if (reset) begin // @[WidthWidget.scala 34:27]
      count <= 1'h0; // @[WidthWidget.scala 34:27]
    end else if (_T) begin // @[WidthWidget.scala 43:24]
      if (last) begin // @[WidthWidget.scala 46:21]
        count <= 1'h0; // @[WidthWidget.scala 47:17]
      end else begin
        count <= count + 1'h1; // @[WidthWidget.scala 44:15]
      end
    end
    if (reset) begin // @[WidthWidget.scala 56:41]
      bundleOut_0_a_bits_data_rdata_written_once <= 1'h0; // @[WidthWidget.scala 56:41]
    end else begin
      bundleOut_0_a_bits_data_rdata_written_once <= _GEN_4;
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 63:35]
      if (bundleOut_0_a_bits_data_masked_enable_0) begin // @[WidthWidget.scala 62:88]
        bundleOut_0_a_bits_data_rdata_0 <= auto_in_a_bits_data;
      end
    end
    if (reset) begin // @[WidthWidget.scala 56:41]
      bundleOut_0_a_bits_mask_rdata_written_once <= 1'h0; // @[WidthWidget.scala 56:41]
    end else begin
      bundleOut_0_a_bits_mask_rdata_written_once <= _GEN_6;
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 63:35]
      if (bundleOut_0_a_bits_mask_masked_enable_0) begin // @[WidthWidget.scala 62:88]
        bundleOut_0_a_bits_mask_rdata_0 <= auto_in_a_bits_mask;
      end
    end
    if (reset) begin // @[WidthWidget.scala 99:26]
      repeat_count <= 1'h0; // @[WidthWidget.scala 99:26]
    end else if (_repeat_T) begin // @[WidthWidget.scala 103:25]
      if (repeat_last) begin // @[WidthWidget.scala 105:21]
        repeat_count <= 1'h0; // @[WidthWidget.scala 105:29]
      end else begin
        repeat_count <= repeat_count + 1'h1; // @[WidthWidget.scala 104:15]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h0 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_0 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h1 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_1 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h2 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_2 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h3 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_3 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h4 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_4 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h5 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_5 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h6 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_6 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h7 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_7 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h8 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_8 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h9 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_9 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'ha == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_10 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'hb == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_11 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'hc == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_12 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'hd == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_13 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'he == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_14 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'hf == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_15 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h10 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_16 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h11 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_17 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h12 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_18 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h13 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_19 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h14 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_20 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h15 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_21 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h16 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_22 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h17 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_23 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h18 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_24 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h19 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_25 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h1a == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_26 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h1b == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_27 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h1c == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_28 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h1d == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_29 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h1e == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_30 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h1f == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_31 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h20 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_32 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h21 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_33 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h22 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_34 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h23 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_35 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h24 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_36 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h25 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_37 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h26 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_38 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h27 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_39 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h28 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_40 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h29 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_41 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h2a == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_42 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h2b == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_43 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h2c == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_44 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h2d == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_45 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h2e == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_46 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h2f == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_47 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h30 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_48 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h31 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_49 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h32 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_50 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h33 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_51 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h34 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_52 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h35 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_53 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h36 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_54 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h37 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_55 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h38 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_56 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h39 == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_57 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h3a == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_58 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h3b == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_59 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h3c == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_60 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h3d == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_61 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h3e == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_62 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 182:28]
      if (6'h3f == auto_in_a_bits_source) begin // @[WidthWidget.scala 183:37]
        repeat_sel_sel_sources_63 <= bundleOut_0_a_bits_mask_bit; // @[WidthWidget.scala 183:37]
      end
    end
    if (repeat_first) begin // @[Reg.scala 16:19]
      if (6'h3f == cated_bits_source) begin // @[Reg.scala 16:23]
        repeat_sel_hold_r <= repeat_sel_sel_sources_63; // @[Reg.scala 16:23]
      end else if (6'h3e == cated_bits_source) begin // @[Reg.scala 16:23]
        repeat_sel_hold_r <= repeat_sel_sel_sources_62; // @[Reg.scala 16:23]
      end else if (6'h3d == cated_bits_source) begin // @[Reg.scala 16:23]
        repeat_sel_hold_r <= repeat_sel_sel_sources_61; // @[Reg.scala 16:23]
      end else begin
        repeat_sel_hold_r <= _GEN_198;
      end
    end
    if (reset) begin // @[WidthWidget.scala 34:27]
      count_1 <= 1'h0; // @[WidthWidget.scala 34:27]
    end else if (_T_1) begin // @[WidthWidget.scala 43:24]
      if (last_1) begin // @[WidthWidget.scala 46:21]
        count_1 <= 1'h0; // @[WidthWidget.scala 47:17]
      end else begin
        count_1 <= count_1 + 1'h1; // @[WidthWidget.scala 44:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bundleOut_0_a_bits_data_rdata_written_once = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bundleOut_0_a_bits_data_rdata_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bundleOut_0_a_bits_mask_rdata_written_once = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bundleOut_0_a_bits_mask_rdata_0 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  repeat_count = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  repeat_sel_sel_sources_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  repeat_sel_sel_sources_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  repeat_sel_sel_sources_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  repeat_sel_sel_sources_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  repeat_sel_sel_sources_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  repeat_sel_sel_sources_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  repeat_sel_sel_sources_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  repeat_sel_sel_sources_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  repeat_sel_sel_sources_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  repeat_sel_sel_sources_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  repeat_sel_sel_sources_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  repeat_sel_sel_sources_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  repeat_sel_sel_sources_12 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  repeat_sel_sel_sources_13 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  repeat_sel_sel_sources_14 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  repeat_sel_sel_sources_15 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  repeat_sel_sel_sources_16 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  repeat_sel_sel_sources_17 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  repeat_sel_sel_sources_18 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  repeat_sel_sel_sources_19 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  repeat_sel_sel_sources_20 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  repeat_sel_sel_sources_21 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  repeat_sel_sel_sources_22 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  repeat_sel_sel_sources_23 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  repeat_sel_sel_sources_24 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  repeat_sel_sel_sources_25 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  repeat_sel_sel_sources_26 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  repeat_sel_sel_sources_27 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  repeat_sel_sel_sources_28 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  repeat_sel_sel_sources_29 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  repeat_sel_sel_sources_30 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  repeat_sel_sel_sources_31 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  repeat_sel_sel_sources_32 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  repeat_sel_sel_sources_33 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  repeat_sel_sel_sources_34 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  repeat_sel_sel_sources_35 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  repeat_sel_sel_sources_36 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  repeat_sel_sel_sources_37 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  repeat_sel_sel_sources_38 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  repeat_sel_sel_sources_39 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  repeat_sel_sel_sources_40 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  repeat_sel_sel_sources_41 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  repeat_sel_sel_sources_42 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  repeat_sel_sel_sources_43 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  repeat_sel_sel_sources_44 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  repeat_sel_sel_sources_45 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  repeat_sel_sel_sources_46 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  repeat_sel_sel_sources_47 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  repeat_sel_sel_sources_48 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  repeat_sel_sel_sources_49 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  repeat_sel_sel_sources_50 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  repeat_sel_sel_sources_51 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  repeat_sel_sel_sources_52 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  repeat_sel_sel_sources_53 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  repeat_sel_sel_sources_54 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  repeat_sel_sel_sources_55 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  repeat_sel_sel_sources_56 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  repeat_sel_sel_sources_57 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  repeat_sel_sel_sources_58 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  repeat_sel_sel_sources_59 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  repeat_sel_sel_sources_60 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  repeat_sel_sel_sources_61 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  repeat_sel_sel_sources_62 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  repeat_sel_sel_sources_63 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  repeat_sel_hold_r = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  count_1 = _RAND_71[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_16(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [12:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_a_bits_corrupt,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [2:0]  io_in_c_bits_size,
  input  [6:0]  io_in_c_bits_source,
  input  [12:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [2:0]  io_in_d_bits_size,
  input  [6:0]  io_in_d_bits_source,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  _source_ok_T_1 = io_in_a_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_7 = io_in_a_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_13 = io_in_a_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_19 = io_in_a_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_25 = io_in_a_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_31 = io_in_a_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_37 = io_in_a_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_43 = io_in_a_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok = _source_ok_T_1 | _source_ok_T_7 | _source_ok_T_13 | _source_ok_T_19 | _source_ok_T_25 |
    _source_ok_T_31 | _source_ok_T_37 | _source_ok_T_43; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46]
  wire [12:0] _GEN_86 = {{7'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  wire [12:0] _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  wire  is_aligned = _is_aligned_T == 13'h0; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  wire  mask_acc = _mask_T | mask_size & mask_nbit; // @[Misc.scala 214:29]
  wire  mask_acc_1 = _mask_T | mask_size & mask_bit; // @[Misc.scala 214:29]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_2 = mask_acc | mask_size_1 & mask_eq_2; // @[Misc.scala 214:29]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_3 = mask_acc | mask_size_1 & mask_eq_3; // @[Misc.scala 214:29]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  wire  mask_acc_4 = mask_acc_1 | mask_size_1 & mask_eq_4; // @[Misc.scala 214:29]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  wire  mask_acc_5 = mask_acc_1 | mask_size_1 & mask_eq_5; // @[Misc.scala 214:29]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_lo = mask_acc_2 | mask_size_2 & mask_eq_6; // @[Misc.scala 214:29]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_lo_hi = mask_acc_2 | mask_size_2 & mask_eq_7; // @[Misc.scala 214:29]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_lo = mask_acc_3 | mask_size_2 & mask_eq_8; // @[Misc.scala 214:29]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_lo_hi_hi = mask_acc_3 | mask_size_2 & mask_eq_9; // @[Misc.scala 214:29]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_lo = mask_acc_4 | mask_size_2 & mask_eq_10; // @[Misc.scala 214:29]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_lo_hi = mask_acc_4 | mask_size_2 & mask_eq_11; // @[Misc.scala 214:29]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_lo = mask_acc_5 | mask_size_2 & mask_eq_12; // @[Misc.scala 214:29]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27]
  wire  mask_hi_hi_hi = mask_acc_5 | mask_size_2 & mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_118 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  wire  _T_180 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire [12:0] _T_183 = io_in_a_bits_address ^ 13'h1000; // @[Parameters.scala 137:31]
  wire [13:0] _T_184 = {1'b0,$signed(_T_183)}; // @[Parameters.scala 137:49]
  wire [13:0] _T_186 = $signed(_T_184) & -14'sh1000; // @[Parameters.scala 137:52]
  wire  _T_187 = $signed(_T_186) == 14'sh0; // @[Parameters.scala 137:67]
  wire  _T_188 = _T_180 & _T_187; // @[Parameters.scala 670:56]
  wire  _T_190 = source_ok & _T_188; // @[Monitor.scala 82:72]
  wire  _T_245 = _source_ok_T_1 & _T_180; // @[Mux.scala 27:72]
  wire  _T_271 = _T_245 & _T_187; // @[Monitor.scala 83:78]
  wire  _T_285 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  wire [7:0] _T_289 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18]
  wire  _T_290 = _T_289 == 8'h0; // @[Monitor.scala 88:31]
  wire  _T_294 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18]
  wire  _T_298 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  wire  _T_469 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  wire  _T_482 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  wire  _T_566 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  wire  _T_570 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  wire  _T_578 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  wire  _T_668 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  wire [7:0] _T_754 = ~mask; // @[Monitor.scala 127:33]
  wire [7:0] _T_755 = io_in_a_bits_mask & _T_754; // @[Monitor.scala 127:31]
  wire  _T_756 = _T_755 == 8'h0; // @[Monitor.scala 127:40]
  wire  _T_760 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  wire  _T_842 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  wire  _T_850 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  wire  _T_932 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  wire  _T_940 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  wire  _T_1022 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  wire  _T_1034 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  wire  _source_ok_T_55 = io_in_d_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_61 = io_in_d_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_67 = io_in_d_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_73 = io_in_d_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_79 = io_in_d_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_85 = io_in_d_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_91 = io_in_d_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_97 = io_in_d_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_1 = _source_ok_T_55 | _source_ok_T_61 | _source_ok_T_67 | _source_ok_T_73 | _source_ok_T_79 |
    _source_ok_T_85 | _source_ok_T_91 | _source_ok_T_97; // @[Parameters.scala 1125:46]
  wire  _T_1038 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  wire  _T_1042 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27]
  wire  _T_1046 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  wire  _T_1050 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15]
  wire  _T_1054 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15]
  wire  _T_1058 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  wire  _T_1069 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  wire  _T_1073 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  wire  _T_1086 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  wire  _T_1106 = _T_1054 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  wire  _T_1115 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  wire  _T_1132 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  wire  _T_1150 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  wire  _source_ok_T_109 = io_in_c_bits_source[6:4] == 3'h0; // @[Parameters.scala 54:32]
  wire  _source_ok_T_115 = io_in_c_bits_source[6:4] == 3'h1; // @[Parameters.scala 54:32]
  wire  _source_ok_T_121 = io_in_c_bits_source[6:4] == 3'h2; // @[Parameters.scala 54:32]
  wire  _source_ok_T_127 = io_in_c_bits_source[6:4] == 3'h3; // @[Parameters.scala 54:32]
  wire  _source_ok_T_133 = io_in_c_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  _source_ok_T_139 = io_in_c_bits_source[6:4] == 3'h5; // @[Parameters.scala 54:32]
  wire  _source_ok_T_145 = io_in_c_bits_source[6:4] == 3'h6; // @[Parameters.scala 54:32]
  wire  _source_ok_T_151 = io_in_c_bits_source[6:4] == 3'h7; // @[Parameters.scala 54:32]
  wire  source_ok_2 = _source_ok_T_109 | _source_ok_T_115 | _source_ok_T_121 | _source_ok_T_127 | _source_ok_T_133 |
    _source_ok_T_139 | _source_ok_T_145 | _source_ok_T_151; // @[Parameters.scala 1125:46]
  wire [12:0] _is_aligned_mask_T_7 = 13'h3f << io_in_c_bits_size; // @[package.scala 234:77]
  wire [5:0] is_aligned_mask_2 = ~_is_aligned_mask_T_7[5:0]; // @[package.scala 234:46]
  wire [12:0] _GEN_87 = {{7'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  wire [12:0] _is_aligned_T_2 = io_in_c_bits_address & _GEN_87; // @[Edges.scala 20:16]
  wire  is_aligned_2 = _is_aligned_T_2 == 13'h0; // @[Edges.scala 20:24]
  wire [12:0] _address_ok_T_5 = io_in_c_bits_address ^ 13'h1000; // @[Parameters.scala 137:31]
  wire [13:0] _address_ok_T_6 = {1'b0,$signed(_address_ok_T_5)}; // @[Parameters.scala 137:49]
  wire [13:0] _address_ok_T_8 = $signed(_address_ok_T_6) & -14'sh1000; // @[Parameters.scala 137:52]
  wire  _address_ok_T_9 = $signed(_address_ok_T_8) == 14'sh0; // @[Parameters.scala 137:67]
  wire  _T_1710 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  wire  _T_1717 = io_in_c_bits_size >= 3'h3; // @[Monitor.scala 245:30]
  wire  _T_1724 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  wire  _T_1732 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  wire  _T_1750 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  wire  _T_1812 = io_in_c_bits_size <= 3'h6; // @[Parameters.scala 92:42]
  wire  _T_1820 = _T_1812 & _address_ok_T_9; // @[Parameters.scala 670:56]
  wire  _T_1822 = source_ok_2 & _T_1820; // @[Monitor.scala 260:78]
  wire  _T_1877 = _source_ok_T_109 & _T_1812; // @[Mux.scala 27:72]
  wire  _T_1903 = _T_1877 & _address_ok_T_9; // @[Monitor.scala 261:78]
  wire  _T_1925 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  wire  _T_2096 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  wire  _T_2106 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  wire  _T_2114 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  wire  _T_2128 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [2:0] size; // @[Monitor.scala 386:22]
  reg [6:0] source; // @[Monitor.scala 387:22]
  reg [12:0] address; // @[Monitor.scala 388:22]
  wire  _T_2150 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  wire  _T_2151 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  wire  _T_2155 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  wire  _T_2159 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  wire  _T_2163 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  wire  _T_2167 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [2:0] size_1; // @[Monitor.scala 537:22]
  reg [6:0] source_1; // @[Monitor.scala 538:22]
  reg  denied; // @[Monitor.scala 540:22]
  wire  _T_2174 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  wire  _T_2175 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  wire  _T_2179 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  wire  _T_2183 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  wire  _T_2187 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  wire  _T_2195 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  wire  _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  wire [2:0] c_first_beats1_decode = is_aligned_mask_2[5:3]; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  reg [2:0] c_first_counter; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1 = c_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  c_first = c_first_counter == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [2:0] size_3; // @[Monitor.scala 514:22]
  reg [6:0] source_3; // @[Monitor.scala 515:22]
  reg [12:0] address_2; // @[Monitor.scala 516:22]
  wire  _T_2226 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  wire  _T_2227 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  wire  _T_2231 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  wire  _T_2235 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  wire  _T_2239 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  wire  _T_2243 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  reg [127:0] inflight; // @[Monitor.scala 611:27]
  reg [511:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [511:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  wire [8:0] _GEN_88 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  wire [9:0] _a_opcode_lookup_T = {{1'd0}, _GEN_88}; // @[Monitor.scala 634:69]
  wire [511:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  wire [511:0] _GEN_89 = {{496'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_89; // @[Monitor.scala 634:97]
  wire [511:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[511:1]}; // @[Monitor.scala 634:152]
  wire [511:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40]
  wire [511:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 638:91]
  wire [511:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[511:1]}; // @[Monitor.scala 638:144]
  wire  _T_2249 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  wire [127:0] _a_set_wo_ready_T = 128'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] a_set_wo_ready = io_in_a_valid & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 648:71 Monitor.scala 649:22]
  wire  _T_2252 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59]
  wire [8:0] _GEN_94 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  wire [9:0] _a_opcodes_set_T = {{1'd0}, _GEN_94}; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm = _a_first_T & a_first_1 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 654:28]
  wire [1026:0] _GEN_95 = {{1023'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  wire [1026:0] _a_opcodes_set_T_1 = _GEN_95 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  wire [3:0] a_sizes_set_interm = _a_first_T & a_first_1 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 Monitor.scala 655:28]
  wire [1026:0] _GEN_97 = {{1023'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  wire [1026:0] _a_sizes_set_T_1 = _GEN_97 << _a_opcodes_set_T; // @[Monitor.scala 657:52]
  wire [127:0] _T_2254 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  wire  _T_2256 = ~_T_2254[0]; // @[Monitor.scala 658:17]
  wire [127:0] a_set = _a_first_T & a_first_1 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 652:72 Monitor.scala 653:28]
  wire [1026:0] _GEN_31 = _a_first_T & a_first_1 ? _a_opcodes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 656:28]
  wire [1026:0] _GEN_32 = _a_first_T & a_first_1 ? _a_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 Monitor.scala 657:28]
  wire  _T_2260 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  wire  _T_2262 = ~_T_1038; // @[Monitor.scala 671:74]
  wire  _T_2263 = io_in_d_valid & d_first_1 & ~_T_1038; // @[Monitor.scala 671:71]
  wire [127:0] _d_clr_wo_ready_T = 128'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] d_clr_wo_ready = io_in_d_valid & d_first_1 & ~_T_1038 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 671:90 Monitor.scala 672:22]
  wire [1038:0] _GEN_99 = {{1023'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  wire [1038:0] _d_opcodes_clr_T_5 = _GEN_99 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  wire [127:0] d_clr = _d_first_T & d_first_1 & _T_2262 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 675:91 Monitor.scala 676:21]
  wire [1038:0] _GEN_35 = _d_first_T & d_first_1 & _T_2262 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 675:91 Monitor.scala 677:21]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  wire  same_cycle_resp = _T_2249 & io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:88]
  wire [127:0] _T_2273 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  wire  _T_2275 = _T_2273[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  wire [2:0] _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38 Monitor.scala 685:38]
  wire [2:0] _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire [2:0] _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39 Monitor.scala 686:39]
  wire  _T_2280 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_2281 = io_in_d_bits_opcode == _GEN_44 | _T_2280; // @[Monitor.scala 685:77]
  wire  _T_2285 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0];
  wire [2:0] _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38 Monitor.scala 689:38]
  wire [2:0] _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire [2:0] _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38 Monitor.scala 690:38]
  wire  _T_2292 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_2293 = io_in_d_bits_opcode == _GEN_60 | _T_2292; // @[Monitor.scala 689:72]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0];
  wire [3:0] _GEN_102 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  wire  _T_2297 = _GEN_102 == a_size_lookup; // @[Monitor.scala 691:36]
  wire  _T_2307 = _T_2260 & a_first_1 & io_in_a_valid & _same_cycle_resp_T_2 & _T_2262; // @[Monitor.scala 694:116]
  wire  _T_2308 = ~io_in_d_ready; // @[Monitor.scala 695:15]
  wire  _T_2309 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  wire  _T_2316 = a_set_wo_ready != d_clr_wo_ready | ~(|a_set_wo_ready); // @[Monitor.scala 699:48]
  wire [127:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  wire [127:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38]
  wire [127:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36]
  wire [511:0] a_opcodes_set = _GEN_31[511:0];
  wire [511:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  wire [511:0] d_opcodes_clr = _GEN_35[511:0];
  wire [511:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62]
  wire [511:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60]
  wire [511:0] a_sizes_set = _GEN_32[511:0];
  wire [511:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  wire [511:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  wire  _T_2325 = ~(|inflight) | plusarg_reader_out == 32'h0 | watchdog < plusarg_reader_out; // @[Monitor.scala 709:47]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  reg [127:0] inflight_1; // @[Monitor.scala 723:35]
  reg [511:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [2:0] c_first_counter_1; // @[Edges.scala 228:27]
  wire [2:0] c_first_counter1_1 = c_first_counter_1 - 3'h1; // @[Edges.scala 229:28]
  wire  c_first_1 = c_first_counter_1 == 3'h0; // @[Edges.scala 230:25]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25]
  wire [511:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42]
  wire [511:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_89; // @[Monitor.scala 747:93]
  wire [511:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[511:1]}; // @[Monitor.scala 747:146]
  wire  _T_2335 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  wire  _T_2336 = io_in_c_valid & c_first_1 & _T_2335; // @[Monitor.scala 756:37]
  wire [127:0] _c_set_wo_ready_T = 128'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  wire [127:0] c_set_wo_ready = io_in_c_valid & c_first_1 & _T_2335 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 756:71 Monitor.scala 757:22]
  wire  _T_2342 = _c_first_T & c_first_1 & _T_2335; // @[Monitor.scala 760:38]
  wire [3:0] _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  wire [3:0] _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 4'h1; // @[Monitor.scala 763:59]
  wire [8:0] _GEN_109 = {io_in_c_bits_source, 2'h0}; // @[Monitor.scala 764:79]
  wire [9:0] _c_opcodes_set_T = {{1'd0}, _GEN_109}; // @[Monitor.scala 764:79]
  wire [3:0] c_sizes_set_interm = _c_first_T & c_first_1 & _T_2335 ? _c_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 760:72 Monitor.scala 763:28]
  wire [1026:0] _GEN_112 = {{1023'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  wire [1026:0] _c_sizes_set_T_1 = _GEN_112 << _c_opcodes_set_T; // @[Monitor.scala 765:52]
  wire [127:0] _T_2343 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  wire  _T_2345 = ~_T_2343[0]; // @[Monitor.scala 766:17]
  wire [127:0] c_set = _c_first_T & c_first_1 & _T_2335 ? _c_set_wo_ready_T : 128'h0; // @[Monitor.scala 760:72 Monitor.scala 761:28]
  wire [1026:0] _GEN_77 = _c_first_T & c_first_1 & _T_2335 ? _c_sizes_set_T_1 : 1027'h0; // @[Monitor.scala 760:72 Monitor.scala 765:28]
  wire  _T_2349 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  wire  _T_2351 = io_in_d_valid & d_first_2 & _T_1038; // @[Monitor.scala 779:71]
  wire [127:0] d_clr_wo_ready_1 = io_in_d_valid & d_first_2 & _T_1038 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 779:89 Monitor.scala 780:22]
  wire [127:0] d_clr_1 = _d_first_T & d_first_2 & _T_1038 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 783:90 Monitor.scala 784:21]
  wire [1038:0] _GEN_80 = _d_first_T & d_first_2 & _T_1038 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 783:90 Monitor.scala 785:21]
  wire  _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1 = _T_2336 & io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:88]
  wire [127:0] _T_2359 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  wire  _T_2361 = _T_2359[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  wire  _T_2365 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0];
  wire  _T_2369 = _GEN_102 == c_size_lookup; // @[Monitor.scala 795:36]
  wire  _T_2378 = _T_2349 & c_first_1 & io_in_c_valid & _same_cycle_resp_T_8 & _T_1038; // @[Monitor.scala 799:116]
  wire  _T_2380 = _T_2308 | io_in_c_ready; // @[Monitor.scala 800:32]
  wire  _T_2384 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  wire  _T_2385 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  wire [127:0] _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  wire [127:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46]
  wire [127:0] _inflight_T_5 = _inflight_T_3 & _inflight_T_4; // @[Monitor.scala 809:44]
  wire [511:0] d_opcodes_clr_1 = _GEN_80[511:0];
  wire [511:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62]
  wire [511:0] c_sizes_set = _GEN_77[511:0];
  wire [511:0] _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  wire [511:0] _inflight_sizes_T_5 = _inflight_sizes_T_3 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  wire  _T_2394 = ~(|inflight_1) | plusarg_reader_1_out == 32'h0 | watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:47]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  reg  inflight_2; // @[Monitor.scala 823:27]
  reg [2:0] d_first_counter_3; // @[Edges.scala 228:27]
  wire [2:0] d_first_counter1_3 = d_first_counter_3 - 3'h1; // @[Edges.scala 229:28]
  wire  d_first_3 = d_first_counter_3 == 3'h0; // @[Edges.scala 230:25]
  wire  _T_2406 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  wire  _T_2407 = _d_first_T & d_first_3 & _T_2406; // @[Monitor.scala 829:38]
  wire  _T_2410 = ~inflight_2; // @[Monitor.scala 831:14]
  wire [1:0] _GEN_84 = _d_first_T & d_first_3 & _T_2406 ? 2'h1 : 2'h0; // @[Monitor.scala 829:72 Monitor.scala 830:13]
  wire  d_set = _GEN_84[0];
  wire  _T_2417 = d_set | inflight_2; // @[Monitor.scala 837:24]
  wire [1:0] _GEN_85 = io_in_e_valid ? 2'h1 : 2'h0; // @[Monitor.scala 835:73 Monitor.scala 836:13]
  wire  e_clr = _GEN_85[0];
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15]
    end
    if (_a_first_T & a_first) begin // @[Monitor.scala 396:32]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15]
    end
    if (_d_first_T & d_first) begin // @[Monitor.scala 549:32]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 3'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      opcode_3 <= io_in_c_bits_opcode; // @[Monitor.scala 525:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      param_3 <= io_in_c_bits_param; // @[Monitor.scala 526:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      size_3 <= io_in_c_bits_size; // @[Monitor.scala 527:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      source_3 <= io_in_c_bits_source; // @[Monitor.scala 528:15]
    end
    if (_c_first_T & c_first) begin // @[Monitor.scala 524:32]
      address_2 <= io_in_c_bits_address; // @[Monitor.scala 529:15]
    end
    if (reset) begin // @[Monitor.scala 611:27]
      inflight <= 128'h0; // @[Monitor.scala 611:27]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14]
    end
    if (reset) begin // @[Monitor.scala 613:35]
      inflight_opcodes <= 512'h0; // @[Monitor.scala 613:35]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22]
    end
    if (reset) begin // @[Monitor.scala 615:33]
      inflight_sizes <= 512'h0; // @[Monitor.scala 615:33]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20]
    end
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin // @[Edges.scala 234:17]
      if (a_first_1) begin // @[Edges.scala 235:21]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_1) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27]
      watchdog <= 32'h0; // @[Monitor.scala 706:27]
    end else if (_a_first_T | _d_first_T) begin // @[Monitor.scala 712:47]
      watchdog <= 32'h0; // @[Monitor.scala 712:58]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14]
    end
    if (reset) begin // @[Monitor.scala 723:35]
      inflight_1 <= 128'h0; // @[Monitor.scala 723:35]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22]
    end
    if (reset) begin // @[Monitor.scala 725:35]
      inflight_sizes_1 <= 512'h0; // @[Monitor.scala 725:35]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      c_first_counter_1 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_c_first_T) begin // @[Edges.scala 234:17]
      if (c_first_1) begin // @[Edges.scala 235:21]
        if (c_first_beats1_opdata) begin // @[Edges.scala 220:14]
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 3'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_2) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27]
    end else if (_c_first_T | _d_first_T) begin // @[Monitor.scala 819:47]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14]
    end
    if (reset) begin // @[Monitor.scala 823:27]
      inflight_2 <= 1'h0; // @[Monitor.scala 823:27]
    end else begin
      inflight_2 <= (inflight_2 | d_set) & ~e_clr; // @[Monitor.scala 842:14]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter_3 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin // @[Edges.scala 234:17]
      if (d_first_3) begin // @[Edges.scala 235:21]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14]
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 3'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_271 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_271 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_285 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_285 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_290 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_290 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_294 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_118 & ~(_T_294 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_271 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_271 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_mask_T | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_mask_T | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_285 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_285 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_469 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_469 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_290 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_290 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_294 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_298 & ~(_T_294 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_188 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_188 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_566 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_566 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_294 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_482 & ~(_T_294 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_566 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_566 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_578 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_566 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_566 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_756 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_668 & ~(_T_756 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_842 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_842 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_760 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_932 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_932 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_850 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_190 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_190 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(source_ok | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(source_ok | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(is_aligned | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(is_aligned | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_1022 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_1022 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_570 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_570 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_294 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & _T_940 & ~(_T_294 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1034 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~(_T_1034 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1042 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1042 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1046 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1046 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1054 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1038 & ~(_T_1054 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1042 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1042 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1069 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1069 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1073 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1073 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1058 & ~(_T_1050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1042 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1042 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1069 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1069 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1073 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1073 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1086 & ~(_T_1106 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(_T_1046 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(_T_1046 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(_T_1050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1115 & ~(_T_1050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(_T_1046 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(_T_1046 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(_T_1106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1132 & ~(_T_1106 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(source_ok_1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(source_ok_1 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(_T_1046 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(_T_1046 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(_T_1050 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_1150 & ~(_T_1050 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_T_1717 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_T_1717 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_T_1724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1710 & ~(_T_1724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_T_1717 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_T_1717 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_T_1724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1732 & ~(_T_1724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1822 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1822 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1903 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1903 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1717 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1717 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel Release carries invalid report param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1750 & ~(_T_1724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1822 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1822 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1903 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1903 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1717 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1717 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1724 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_1925 & ~(_T_1724 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(_T_2106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2096 & ~(_T_2106 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(_T_2106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2114 & ~(_T_2106 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(_address_ok_T_9 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(_address_ok_T_9 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(source_ok_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(source_ok_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(is_aligned_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(is_aligned_2 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(_T_2106 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel HintAck carries invalid param (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_c_valid & _T_2128 & ~(_T_2106 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2151 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2151 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2155 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2155 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2159 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2159 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2163 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2163 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2150 & ~(_T_2167 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2150 & ~(_T_2167 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2175 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2175 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2179 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2179 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2183 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2183 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2187 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2187 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & ~(_T_2195 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & ~(_T_2195 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2227 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2227 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2231 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel param changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2231 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2235 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel size changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2235 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2239 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel source changed within multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2239 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2226 & ~(_T_2243 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel address changed with multibeat operation (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2226 & ~(_T_2243 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2252 & ~(_T_2256 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2252 & ~(_T_2256 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & ~(_T_2275 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & ~(_T_2275 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & same_cycle_resp & ~(_T_2281 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & same_cycle_resp & ~(_T_2281 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & same_cycle_resp & ~(_T_2285 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & same_cycle_resp & ~(_T_2285 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & ~same_cycle_resp & ~(_T_2293 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & ~same_cycle_resp & ~(_T_2293 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2263 & ~same_cycle_resp & ~(_T_2297 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2263 & ~same_cycle_resp & ~(_T_2297 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2307 & ~(_T_2309 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2307 & ~(_T_2309 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2316 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2316 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2325 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2325 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2342 & ~(_T_2345 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' channel re-used a source ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2342 & ~(_T_2345 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2351 & ~(_T_2361 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2351 & ~(_T_2361 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2351 & same_cycle_resp_1 & ~(_T_2365 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2351 & same_cycle_resp_1 & ~(_T_2365 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2351 & ~same_cycle_resp_1 & ~(_T_2369 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2351 & ~same_cycle_resp_1 & ~(_T_2369 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2378 & ~(_T_2380 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2378 & ~(_T_2380 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2384 & ~(_T_2385 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2384 & ~(_T_2385 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_2394 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_2394 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2407 & ~(_T_2410 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel re-used a sink ID (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2407 & ~(_T_2410 | reset)) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & ~(_T_2417 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChipLinkBridge.scala:154:32)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & ~(_T_2417 | reset)) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  denied = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  c_first_counter = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  opcode_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  param_3 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  size_3 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  source_3 = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  address_2 = _RAND_17[12:0];
  _RAND_18 = {4{`RANDOM}};
  inflight = _RAND_18[127:0];
  _RAND_19 = {16{`RANDOM}};
  inflight_opcodes = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  inflight_sizes = _RAND_20[511:0];
  _RAND_21 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  watchdog = _RAND_23[31:0];
  _RAND_24 = {4{`RANDOM}};
  inflight_1 = _RAND_24[127:0];
  _RAND_25 = {16{`RANDOM}};
  inflight_sizes_1 = _RAND_25[511:0];
  _RAND_26 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  watchdog_1 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inflight_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_30[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_4(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [12:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [12:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output        io_deq_bits_corrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_param; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [6:0] saved_source; // @[Repeater.scala 20:18]
  reg [12:0] saved_address; // @[Repeater.scala 20:18]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18]
  reg  saved_corrupt; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 28:38 Repeater.scala 28:45 Repeater.scala 19:21]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; // @[Repeater.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin // @[Repeater.scala 29:38]
      full <= 1'h0; // @[Repeater.scala 29:45]
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_param <= io_enq_bits_param; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_corrupt <= io_enq_bits_corrupt; // @[Repeater.scala 28:62]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  saved_mask = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  saved_corrupt = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_5(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [12:0] io_enq_bits_address,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [12:0] io_deq_bits_address
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_param; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [6:0] saved_source; // @[Repeater.scala 20:18]
  reg [12:0] saved_address; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 28:38 Repeater.scala 28:45 Repeater.scala 19:21]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin // @[Repeater.scala 29:38]
      full <= 1'h0; // @[Repeater.scala 29:45]
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_param <= io_enq_bits_param; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[12:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLWidthWidget_2(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [12:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input         auto_in_a_bits_corrupt,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [2:0]  auto_in_c_bits_size,
  input  [6:0]  auto_in_c_bits_source,
  input  [12:0] auto_in_c_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output        auto_in_d_bits_corrupt,
  input         auto_in_e_valid,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [2:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [12:0] auto_out_a_bits_address,
  output [3:0]  auto_out_a_bits_mask,
  output        auto_out_a_bits_corrupt,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [2:0]  auto_out_c_bits_size,
  output [6:0]  auto_out_c_bits_source,
  output [12:0] auto_out_c_bits_address,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [2:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input         auto_out_d_bits_corrupt,
  output        auto_out_e_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [12:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [12:0] monitor_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [6:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_valid; // @[Nodes.scala 24:25]
  wire  repeated_repeater_clock; // @[Repeater.scala 35:26]
  wire  repeated_repeater_reset; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_repeat; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_param; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_size; // @[Repeater.scala 35:26]
  wire [6:0] repeated_repeater_io_enq_bits_source; // @[Repeater.scala 35:26]
  wire [12:0] repeated_repeater_io_enq_bits_address; // @[Repeater.scala 35:26]
  wire [7:0] repeated_repeater_io_enq_bits_mask; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_bits_corrupt; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_param; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_size; // @[Repeater.scala 35:26]
  wire [6:0] repeated_repeater_io_deq_bits_source; // @[Repeater.scala 35:26]
  wire [12:0] repeated_repeater_io_deq_bits_address; // @[Repeater.scala 35:26]
  wire [7:0] repeated_repeater_io_deq_bits_mask; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_bits_corrupt; // @[Repeater.scala 35:26]
  wire  repeated_repeater_1_clock; // @[Repeater.scala 35:26]
  wire  repeated_repeater_1_reset; // @[Repeater.scala 35:26]
  wire  repeated_repeater_1_io_repeat; // @[Repeater.scala 35:26]
  wire  repeated_repeater_1_io_enq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_1_io_enq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_1_io_enq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_1_io_enq_bits_param; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_1_io_enq_bits_size; // @[Repeater.scala 35:26]
  wire [6:0] repeated_repeater_1_io_enq_bits_source; // @[Repeater.scala 35:26]
  wire [12:0] repeated_repeater_1_io_enq_bits_address; // @[Repeater.scala 35:26]
  wire  repeated_repeater_1_io_deq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_1_io_deq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_1_io_deq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_1_io_deq_bits_param; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_1_io_deq_bits_size; // @[Repeater.scala 35:26]
  wire [6:0] repeated_repeater_1_io_deq_bits_source; // @[Repeater.scala 35:26]
  wire [12:0] repeated_repeater_1_io_deq_bits_address; // @[Repeater.scala 35:26]
  wire [2:0] cated_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  repeat_hasData = ~cated_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] cated_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire [9:0] _repeat_limit_T_1 = 10'h7 << cated_bits_size; // @[package.scala 234:77]
  wire [2:0] _repeat_limit_T_3 = ~_repeat_limit_T_1[2:0]; // @[package.scala 234:46]
  wire  repeat_limit = _repeat_limit_T_3[2]; // @[WidthWidget.scala 97:47]
  reg  repeat_count; // @[WidthWidget.scala 99:26]
  wire  repeat_last = repeat_count == repeat_limit | ~repeat_hasData; // @[WidthWidget.scala 101:35]
  wire  cated_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  _repeat_T = auto_out_a_ready & cated_valid; // @[Decoupled.scala 40:37]
  wire [12:0] cated_bits_address = repeated_repeater_io_deq_bits_address; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  repeat_sel = cated_bits_address[2]; // @[WidthWidget.scala 110:39]
  wire  repeat_index = repeat_sel | repeat_count; // @[WidthWidget.scala 120:24]
  wire [7:0] cated_bits_mask = repeated_repeater_io_deq_bits_mask; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire [3:0] repeat_bundleOut_0_a_bits_mask_mux_0 = cated_bits_mask[3:0]; // @[WidthWidget.scala 122:55]
  wire [3:0] repeat_bundleOut_0_a_bits_mask_mux_1 = cated_bits_mask[7:4]; // @[WidthWidget.scala 122:55]
  wire  hasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [9:0] _limit_T_1 = 10'h7 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [2:0] _limit_T_3 = ~_limit_T_1[2:0]; // @[package.scala 234:46]
  wire  limit = _limit_T_3[2]; // @[WidthWidget.scala 32:47]
  reg  count; // @[WidthWidget.scala 34:27]
  wire  last = count == limit | ~hasData; // @[WidthWidget.scala 36:36]
  reg  corrupt_reg; // @[WidthWidget.scala 39:32]
  wire  corrupt_out = auto_out_d_bits_corrupt | corrupt_reg; // @[WidthWidget.scala 41:36]
  wire  bundleOut_0_d_ready = auto_in_d_ready | ~last; // @[WidthWidget.scala 70:29]
  wire  _T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  wire [2:0] cated_1_bits_opcode = repeated_repeater_1_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  repeat_hasData_1 = cated_1_bits_opcode[0]; // @[Edges.scala 101:36]
  wire [2:0] cated_1_bits_size = repeated_repeater_1_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire [9:0] _repeat_limit_T_5 = 10'h7 << cated_1_bits_size; // @[package.scala 234:77]
  wire [2:0] _repeat_limit_T_7 = ~_repeat_limit_T_5[2:0]; // @[package.scala 234:46]
  wire  repeat_limit_1 = _repeat_limit_T_7[2]; // @[WidthWidget.scala 97:47]
  reg  repeat_count_1; // @[WidthWidget.scala 99:26]
  wire  repeat_last_1 = repeat_count_1 == repeat_limit_1 | ~repeat_hasData_1; // @[WidthWidget.scala 101:35]
  wire  cated_1_valid = repeated_repeater_1_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  wire  _repeat_T_2 = auto_out_c_ready & cated_1_valid; // @[Decoupled.scala 40:37]
  TLMonitor_16 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_c_ready(monitor_io_in_c_ready),
    .io_in_c_valid(monitor_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_io_in_c_bits_address),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),
    .io_in_e_valid(monitor_io_in_e_valid)
  );
  Repeater_4 repeated_repeater ( // @[Repeater.scala 35:26]
    .clock(repeated_repeater_clock),
    .reset(repeated_repeater_reset),
    .io_repeat(repeated_repeater_io_repeat),
    .io_enq_ready(repeated_repeater_io_enq_ready),
    .io_enq_valid(repeated_repeater_io_enq_valid),
    .io_enq_bits_opcode(repeated_repeater_io_enq_bits_opcode),
    .io_enq_bits_param(repeated_repeater_io_enq_bits_param),
    .io_enq_bits_size(repeated_repeater_io_enq_bits_size),
    .io_enq_bits_source(repeated_repeater_io_enq_bits_source),
    .io_enq_bits_address(repeated_repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeated_repeater_io_enq_bits_mask),
    .io_enq_bits_corrupt(repeated_repeater_io_enq_bits_corrupt),
    .io_deq_ready(repeated_repeater_io_deq_ready),
    .io_deq_valid(repeated_repeater_io_deq_valid),
    .io_deq_bits_opcode(repeated_repeater_io_deq_bits_opcode),
    .io_deq_bits_param(repeated_repeater_io_deq_bits_param),
    .io_deq_bits_size(repeated_repeater_io_deq_bits_size),
    .io_deq_bits_source(repeated_repeater_io_deq_bits_source),
    .io_deq_bits_address(repeated_repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeated_repeater_io_deq_bits_mask),
    .io_deq_bits_corrupt(repeated_repeater_io_deq_bits_corrupt)
  );
  Repeater_5 repeated_repeater_1 ( // @[Repeater.scala 35:26]
    .clock(repeated_repeater_1_clock),
    .reset(repeated_repeater_1_reset),
    .io_repeat(repeated_repeater_1_io_repeat),
    .io_enq_ready(repeated_repeater_1_io_enq_ready),
    .io_enq_valid(repeated_repeater_1_io_enq_valid),
    .io_enq_bits_opcode(repeated_repeater_1_io_enq_bits_opcode),
    .io_enq_bits_param(repeated_repeater_1_io_enq_bits_param),
    .io_enq_bits_size(repeated_repeater_1_io_enq_bits_size),
    .io_enq_bits_source(repeated_repeater_1_io_enq_bits_source),
    .io_enq_bits_address(repeated_repeater_1_io_enq_bits_address),
    .io_deq_ready(repeated_repeater_1_io_deq_ready),
    .io_deq_valid(repeated_repeater_1_io_deq_valid),
    .io_deq_bits_opcode(repeated_repeater_1_io_deq_bits_opcode),
    .io_deq_bits_param(repeated_repeater_1_io_deq_bits_param),
    .io_deq_bits_size(repeated_repeater_1_io_deq_bits_size),
    .io_deq_bits_source(repeated_repeater_1_io_deq_bits_source),
    .io_deq_bits_address(repeated_repeater_1_io_deq_bits_address)
  );
  assign auto_in_a_ready = repeated_repeater_io_enq_ready; // @[Nodes.scala 1210:84 Repeater.scala 37:21]
  assign auto_in_c_ready = repeated_repeater_1_io_enq_ready; // @[Nodes.scala 1210:84 Repeater.scala 37:21]
  assign auto_in_d_valid = auto_out_d_valid & last; // @[WidthWidget.scala 71:29]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt | corrupt_reg; // @[WidthWidget.scala 41:36]
  assign auto_out_a_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_param = repeated_repeater_io_deq_bits_param; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_source = repeated_repeater_io_deq_bits_source; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_address = repeated_repeater_io_deq_bits_address; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_a_bits_mask = repeat_index ? repeat_bundleOut_0_a_bits_mask_mux_1 :
    repeat_bundleOut_0_a_bits_mask_mux_0; // @[WidthWidget.scala 134:53 WidthWidget.scala 134:53]
  assign auto_out_a_bits_corrupt = repeated_repeater_io_deq_bits_corrupt; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_c_valid = repeated_repeater_1_io_deq_valid; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_c_bits_opcode = repeated_repeater_1_io_deq_bits_opcode; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_c_bits_param = repeated_repeater_1_io_deq_bits_param; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_c_bits_size = repeated_repeater_1_io_deq_bits_size; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_c_bits_source = repeated_repeater_1_io_deq_bits_source; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_c_bits_address = repeated_repeater_1_io_deq_bits_address; // @[WidthWidget.scala 155:25 WidthWidget.scala 156:15]
  assign auto_out_d_ready = auto_in_d_ready | ~last; // @[WidthWidget.scala 70:29]
  assign auto_out_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = repeated_repeater_io_enq_ready; // @[Nodes.scala 1210:84 Repeater.scala 37:21]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_ready = repeated_repeater_1_io_enq_ready; // @[Nodes.scala 1210:84 Repeater.scala 37:21]
  assign monitor_io_in_c_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_c_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign monitor_io_in_d_valid = auto_out_d_valid & last; // @[WidthWidget.scala 71:29]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt | corrupt_reg; // @[WidthWidget.scala 41:36]
  assign monitor_io_in_e_valid = auto_in_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_clock = clock;
  assign repeated_repeater_reset = reset;
  assign repeated_repeater_io_repeat = ~repeat_last; // @[WidthWidget.scala 142:7]
  assign repeated_repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign repeated_repeater_1_clock = clock;
  assign repeated_repeater_1_reset = reset;
  assign repeated_repeater_1_io_repeat = ~repeat_last_1; // @[WidthWidget.scala 142:7]
  assign repeated_repeater_1_io_enq_valid = auto_in_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_1_io_enq_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_1_io_enq_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_1_io_enq_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_1_io_enq_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_1_io_enq_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_1_io_deq_ready = auto_out_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  always @(posedge clock) begin
    if (reset) begin // @[WidthWidget.scala 99:26]
      repeat_count <= 1'h0; // @[WidthWidget.scala 99:26]
    end else if (_repeat_T) begin // @[WidthWidget.scala 103:25]
      if (repeat_last) begin // @[WidthWidget.scala 105:21]
        repeat_count <= 1'h0; // @[WidthWidget.scala 105:29]
      end else begin
        repeat_count <= repeat_count + 1'h1; // @[WidthWidget.scala 104:15]
      end
    end
    if (reset) begin // @[WidthWidget.scala 34:27]
      count <= 1'h0; // @[WidthWidget.scala 34:27]
    end else if (_T) begin // @[WidthWidget.scala 43:24]
      if (last) begin // @[WidthWidget.scala 46:21]
        count <= 1'h0; // @[WidthWidget.scala 47:17]
      end else begin
        count <= count + 1'h1; // @[WidthWidget.scala 44:15]
      end
    end
    if (reset) begin // @[WidthWidget.scala 39:32]
      corrupt_reg <= 1'h0; // @[WidthWidget.scala 39:32]
    end else if (_T) begin // @[WidthWidget.scala 43:24]
      if (last) begin // @[WidthWidget.scala 46:21]
        corrupt_reg <= 1'h0; // @[WidthWidget.scala 48:23]
      end else begin
        corrupt_reg <= corrupt_out; // @[WidthWidget.scala 45:21]
      end
    end
    if (reset) begin // @[WidthWidget.scala 99:26]
      repeat_count_1 <= 1'h0; // @[WidthWidget.scala 99:26]
    end else if (_repeat_T_2) begin // @[WidthWidget.scala 103:25]
      if (repeat_last_1) begin // @[WidthWidget.scala 105:21]
        repeat_count_1 <= 1'h0; // @[WidthWidget.scala 105:29]
      end else begin
        repeat_count_1 <= repeat_count_1 + 1'h1; // @[WidthWidget.scala 104:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  repeat_count = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  corrupt_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  repeat_count_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ChipLinkMaster(
  input         clock,
  input         reset,
  output        slave_0_awready,
  input         slave_0_awvalid,
  input  [3:0]  slave_0_awid,
  input  [31:0] slave_0_awaddr,
  input  [7:0]  slave_0_awlen,
  input  [2:0]  slave_0_awsize,
  input  [1:0]  slave_0_awburst,
  output        slave_0_wready,
  input         slave_0_wvalid,
  input  [63:0] slave_0_wdata,
  input  [7:0]  slave_0_wstrb,
  input         slave_0_wlast,
  input         slave_0_bready,
  output        slave_0_bvalid,
  output [3:0]  slave_0_bid,
  output [1:0]  slave_0_bresp,
  output        slave_0_arready,
  input         slave_0_arvalid,
  input  [3:0]  slave_0_arid,
  input  [31:0] slave_0_araddr,
  input  [7:0]  slave_0_arlen,
  input  [2:0]  slave_0_arsize,
  input  [1:0]  slave_0_arburst,
  input         slave_0_rready,
  output        slave_0_rvalid,
  output [3:0]  slave_0_rid,
  output [63:0] slave_0_rdata,
  output [1:0]  slave_0_rresp,
  output        slave_0_rlast,
  input         master_mem_0_awready,
  output        master_mem_0_awvalid,
  output [3:0]  master_mem_0_awid,
  output [31:0] master_mem_0_awaddr,
  output [7:0]  master_mem_0_awlen,
  output [2:0]  master_mem_0_awsize,
  output [1:0]  master_mem_0_awburst,
  input         master_mem_0_wready,
  output        master_mem_0_wvalid,
  output [63:0] master_mem_0_wdata,
  output [7:0]  master_mem_0_wstrb,
  output        master_mem_0_wlast,
  output        master_mem_0_bready,
  input         master_mem_0_bvalid,
  input  [3:0]  master_mem_0_bid,
  input  [1:0]  master_mem_0_bresp,
  input         master_mem_0_arready,
  output        master_mem_0_arvalid,
  output [3:0]  master_mem_0_arid,
  output [31:0] master_mem_0_araddr,
  output [7:0]  master_mem_0_arlen,
  output [2:0]  master_mem_0_arsize,
  output [1:0]  master_mem_0_arburst,
  output        master_mem_0_rready,
  input         master_mem_0_rvalid,
  input  [3:0]  master_mem_0_rid,
  input  [63:0] master_mem_0_rdata,
  input  [1:0]  master_mem_0_rresp,
  input         master_mem_0_rlast,
  output        fpga_io_c2b_clk,
  output        fpga_io_c2b_rst,
  output        fpga_io_c2b_send,
  output [7:0]  fpga_io_c2b_data,
  input         fpga_io_b2c_clk,
  input         fpga_io_b2c_rst,
  input         fpga_io_b2c_send,
  input  [7:0]  fpga_io_b2c_data
);
  wire  xbar_clock; // @[Xbar.scala 142:26]
  wire  xbar_reset; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_a_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_a_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_in_a_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_in_a_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_in_a_bits_size; // @[Xbar.scala 142:26]
  wire [6:0] xbar_auto_in_a_bits_source; // @[Xbar.scala 142:26]
  wire [31:0] xbar_auto_in_a_bits_address; // @[Xbar.scala 142:26]
  wire [7:0] xbar_auto_in_a_bits_mask; // @[Xbar.scala 142:26]
  wire [63:0] xbar_auto_in_a_bits_data; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_a_bits_corrupt; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_c_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_c_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_in_c_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_in_c_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_in_c_bits_size; // @[Xbar.scala 142:26]
  wire [6:0] xbar_auto_in_c_bits_source; // @[Xbar.scala 142:26]
  wire [31:0] xbar_auto_in_c_bits_address; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_d_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_d_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_in_d_bits_opcode; // @[Xbar.scala 142:26]
  wire [1:0] xbar_auto_in_d_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_in_d_bits_size; // @[Xbar.scala 142:26]
  wire [6:0] xbar_auto_in_d_bits_source; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_d_bits_denied; // @[Xbar.scala 142:26]
  wire [63:0] xbar_auto_in_d_bits_data; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_d_bits_corrupt; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_e_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_e_valid; // @[Xbar.scala 142:26]
  wire  xbar_auto_in_e_bits_sink; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_a_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_a_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_1_a_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_1_a_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_1_a_bits_size; // @[Xbar.scala 142:26]
  wire [6:0] xbar_auto_out_1_a_bits_source; // @[Xbar.scala 142:26]
  wire [12:0] xbar_auto_out_1_a_bits_address; // @[Xbar.scala 142:26]
  wire [7:0] xbar_auto_out_1_a_bits_mask; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_a_bits_corrupt; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_c_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_c_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_1_c_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_1_c_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_1_c_bits_size; // @[Xbar.scala 142:26]
  wire [6:0] xbar_auto_out_1_c_bits_source; // @[Xbar.scala 142:26]
  wire [12:0] xbar_auto_out_1_c_bits_address; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_d_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_d_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_1_d_bits_opcode; // @[Xbar.scala 142:26]
  wire [1:0] xbar_auto_out_1_d_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_1_d_bits_size; // @[Xbar.scala 142:26]
  wire [6:0] xbar_auto_out_1_d_bits_source; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_d_bits_denied; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_d_bits_corrupt; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_1_e_valid; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_0_a_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_0_a_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_0_a_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_0_a_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_0_a_bits_size; // @[Xbar.scala 142:26]
  wire [6:0] xbar_auto_out_0_a_bits_source; // @[Xbar.scala 142:26]
  wire [31:0] xbar_auto_out_0_a_bits_address; // @[Xbar.scala 142:26]
  wire [7:0] xbar_auto_out_0_a_bits_mask; // @[Xbar.scala 142:26]
  wire [63:0] xbar_auto_out_0_a_bits_data; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_0_a_bits_corrupt; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_0_d_ready; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_0_d_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_0_d_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_auto_out_0_d_bits_size; // @[Xbar.scala 142:26]
  wire [6:0] xbar_auto_out_0_d_bits_source; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_0_d_bits_denied; // @[Xbar.scala 142:26]
  wire [63:0] xbar_auto_out_0_d_bits_data; // @[Xbar.scala 142:26]
  wire  xbar_auto_out_0_d_bits_corrupt; // @[Xbar.scala 142:26]
  wire  xbar_1_clock; // @[Xbar.scala 142:26]
  wire  xbar_1_reset; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_in_a_ready; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_in_a_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_in_a_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_in_a_bits_size; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_in_a_bits_source; // @[Xbar.scala 142:26]
  wire [31:0] xbar_1_auto_in_a_bits_address; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_in_a_bits_mask; // @[Xbar.scala 142:26]
  wire [31:0] xbar_1_auto_in_a_bits_data; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_in_d_ready; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_in_d_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_in_d_bits_opcode; // @[Xbar.scala 142:26]
  wire [1:0] xbar_1_auto_in_d_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_in_d_bits_size; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_in_d_bits_source; // @[Xbar.scala 142:26]
  wire [5:0] xbar_1_auto_in_d_bits_sink; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_in_d_bits_denied; // @[Xbar.scala 142:26]
  wire [31:0] xbar_1_auto_in_d_bits_data; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_in_d_bits_corrupt; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_1_a_ready; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_1_a_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_out_1_a_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_out_1_a_bits_size; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_out_1_a_bits_source; // @[Xbar.scala 142:26]
  wire [12:0] xbar_1_auto_out_1_a_bits_address; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_out_1_a_bits_mask; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_1_d_ready; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_1_d_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_out_1_d_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_out_1_d_bits_size; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_out_1_d_bits_source; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_1_d_bits_denied; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_1_d_bits_corrupt; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_0_a_ready; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_0_a_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_out_0_a_bits_opcode; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_out_0_a_bits_size; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_out_0_a_bits_source; // @[Xbar.scala 142:26]
  wire [31:0] xbar_1_auto_out_0_a_bits_address; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_out_0_a_bits_mask; // @[Xbar.scala 142:26]
  wire [31:0] xbar_1_auto_out_0_a_bits_data; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_0_d_ready; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_0_d_valid; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_out_0_d_bits_opcode; // @[Xbar.scala 142:26]
  wire [1:0] xbar_1_auto_out_0_d_bits_param; // @[Xbar.scala 142:26]
  wire [2:0] xbar_1_auto_out_0_d_bits_size; // @[Xbar.scala 142:26]
  wire [3:0] xbar_1_auto_out_0_d_bits_source; // @[Xbar.scala 142:26]
  wire [4:0] xbar_1_auto_out_0_d_bits_sink; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_0_d_bits_denied; // @[Xbar.scala 142:26]
  wire [31:0] xbar_1_auto_out_0_d_bits_data; // @[Xbar.scala 142:26]
  wire  xbar_1_auto_out_0_d_bits_corrupt; // @[Xbar.scala 142:26]
  wire  ferr_clock; // @[ChipLinkBridge.scala 31:24]
  wire  ferr_reset; // @[ChipLinkBridge.scala 31:24]
  wire  ferr_auto_in_a_ready; // @[ChipLinkBridge.scala 31:24]
  wire  ferr_auto_in_a_valid; // @[ChipLinkBridge.scala 31:24]
  wire [2:0] ferr_auto_in_a_bits_opcode; // @[ChipLinkBridge.scala 31:24]
  wire [2:0] ferr_auto_in_a_bits_size; // @[ChipLinkBridge.scala 31:24]
  wire [3:0] ferr_auto_in_a_bits_source; // @[ChipLinkBridge.scala 31:24]
  wire [12:0] ferr_auto_in_a_bits_address; // @[ChipLinkBridge.scala 31:24]
  wire [3:0] ferr_auto_in_a_bits_mask; // @[ChipLinkBridge.scala 31:24]
  wire  ferr_auto_in_d_ready; // @[ChipLinkBridge.scala 31:24]
  wire  ferr_auto_in_d_valid; // @[ChipLinkBridge.scala 31:24]
  wire [2:0] ferr_auto_in_d_bits_opcode; // @[ChipLinkBridge.scala 31:24]
  wire [2:0] ferr_auto_in_d_bits_size; // @[ChipLinkBridge.scala 31:24]
  wire [3:0] ferr_auto_in_d_bits_source; // @[ChipLinkBridge.scala 31:24]
  wire  ferr_auto_in_d_bits_denied; // @[ChipLinkBridge.scala 31:24]
  wire  ferr_auto_in_d_bits_corrupt; // @[ChipLinkBridge.scala 31:24]
  wire  chiplink_clock; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_reset; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_a_ready; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_a_valid; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_mbypass_out_a_bits_opcode; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_mbypass_out_a_bits_param; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_mbypass_out_a_bits_size; // @[ChipLinkBridge.scala 39:28]
  wire [5:0] chiplink_auto_mbypass_out_a_bits_source; // @[ChipLinkBridge.scala 39:28]
  wire [31:0] chiplink_auto_mbypass_out_a_bits_address; // @[ChipLinkBridge.scala 39:28]
  wire [3:0] chiplink_auto_mbypass_out_a_bits_mask; // @[ChipLinkBridge.scala 39:28]
  wire [31:0] chiplink_auto_mbypass_out_a_bits_data; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_c_ready; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_c_valid; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_mbypass_out_c_bits_opcode; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_mbypass_out_c_bits_param; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_mbypass_out_c_bits_size; // @[ChipLinkBridge.scala 39:28]
  wire [5:0] chiplink_auto_mbypass_out_c_bits_source; // @[ChipLinkBridge.scala 39:28]
  wire [31:0] chiplink_auto_mbypass_out_c_bits_address; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_d_ready; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_d_valid; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_mbypass_out_d_bits_opcode; // @[ChipLinkBridge.scala 39:28]
  wire [1:0] chiplink_auto_mbypass_out_d_bits_param; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_mbypass_out_d_bits_size; // @[ChipLinkBridge.scala 39:28]
  wire [5:0] chiplink_auto_mbypass_out_d_bits_source; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_d_bits_denied; // @[ChipLinkBridge.scala 39:28]
  wire [31:0] chiplink_auto_mbypass_out_d_bits_data; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_d_bits_corrupt; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_e_ready; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_e_valid; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_mbypass_out_e_bits_sink; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_sbypass_node_in_in_a_ready; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_sbypass_node_in_in_a_valid; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_sbypass_node_in_in_a_bits_opcode; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_sbypass_node_in_in_a_bits_size; // @[ChipLinkBridge.scala 39:28]
  wire [3:0] chiplink_auto_sbypass_node_in_in_a_bits_source; // @[ChipLinkBridge.scala 39:28]
  wire [31:0] chiplink_auto_sbypass_node_in_in_a_bits_address; // @[ChipLinkBridge.scala 39:28]
  wire [3:0] chiplink_auto_sbypass_node_in_in_a_bits_mask; // @[ChipLinkBridge.scala 39:28]
  wire [31:0] chiplink_auto_sbypass_node_in_in_a_bits_data; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_sbypass_node_in_in_d_ready; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_sbypass_node_in_in_d_valid; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_sbypass_node_in_in_d_bits_opcode; // @[ChipLinkBridge.scala 39:28]
  wire [1:0] chiplink_auto_sbypass_node_in_in_d_bits_param; // @[ChipLinkBridge.scala 39:28]
  wire [2:0] chiplink_auto_sbypass_node_in_in_d_bits_size; // @[ChipLinkBridge.scala 39:28]
  wire [3:0] chiplink_auto_sbypass_node_in_in_d_bits_source; // @[ChipLinkBridge.scala 39:28]
  wire [4:0] chiplink_auto_sbypass_node_in_in_d_bits_sink; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_sbypass_node_in_in_d_bits_denied; // @[ChipLinkBridge.scala 39:28]
  wire [31:0] chiplink_auto_sbypass_node_in_in_d_bits_data; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_sbypass_node_in_in_d_bits_corrupt; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_io_out_c2b_clk; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_io_out_c2b_rst; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_io_out_c2b_send; // @[ChipLinkBridge.scala 39:28]
  wire [7:0] chiplink_auto_io_out_c2b_data; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_io_out_b2c_clk; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_io_out_b2c_rst; // @[ChipLinkBridge.scala 39:28]
  wire  chiplink_auto_io_out_b2c_send; // @[ChipLinkBridge.scala 39:28]
  wire [7:0] chiplink_auto_io_out_b2c_data; // @[ChipLinkBridge.scala 39:28]
  wire  fixer_clock; // @[FIFOFixer.scala 144:27]
  wire  fixer_reset; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_in_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_in_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [1:0] fixer_auto_in_d_bits_param; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_in_d_bits_sink; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_in_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_out_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_out_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [1:0] fixer_auto_out_d_bits_param; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_out_d_bits_sink; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_out_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  widget_clock; // @[WidthWidget.scala 219:28]
  wire  widget_reset; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_a_ready; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_a_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_in_a_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[WidthWidget.scala 219:28]
  wire [3:0] widget_auto_in_a_bits_source; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_auto_in_a_bits_address; // @[WidthWidget.scala 219:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[WidthWidget.scala 219:28]
  wire [63:0] widget_auto_in_a_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_d_ready; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_d_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_in_d_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_in_d_bits_size; // @[WidthWidget.scala 219:28]
  wire [3:0] widget_auto_in_d_bits_source; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_d_bits_denied; // @[WidthWidget.scala 219:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_d_bits_corrupt; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_a_ready; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_a_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_out_a_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[WidthWidget.scala 219:28]
  wire [3:0] widget_auto_out_a_bits_source; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_auto_out_a_bits_address; // @[WidthWidget.scala 219:28]
  wire [3:0] widget_auto_out_a_bits_mask; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_auto_out_a_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_d_ready; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_d_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_out_d_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [1:0] widget_auto_out_d_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[WidthWidget.scala 219:28]
  wire [3:0] widget_auto_out_d_bits_source; // @[WidthWidget.scala 219:28]
  wire [5:0] widget_auto_out_d_bits_sink; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_d_bits_denied; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_auto_out_d_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_d_bits_corrupt; // @[WidthWidget.scala 219:28]
  wire  axi42tl_clock; // @[ToTL.scala 216:29]
  wire  axi42tl_reset; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_awready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_awvalid; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_awid; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_in_awaddr; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_awlen; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_awsize; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_wready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_wvalid; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_in_wdata; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_wstrb; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_wlast; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_bready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_bvalid; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_bid; // @[ToTL.scala 216:29]
  wire [1:0] axi42tl_auto_in_bresp; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_arready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_arvalid; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_arid; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_in_araddr; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_arlen; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_arsize; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_rready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_rvalid; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_rid; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_in_rdata; // @[ToTL.scala 216:29]
  wire [1:0] axi42tl_auto_in_rresp; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_rlast; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_valid; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_out_a_bits_opcode; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_out_a_bits_size; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_out_a_bits_source; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_out_a_bits_address; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_out_a_bits_mask; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_out_a_bits_data; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_valid; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_out_d_bits_opcode; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_out_d_bits_size; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_out_d_bits_source; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_bits_denied; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_out_d_bits_data; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_bits_corrupt; // @[ToTL.scala 216:29]
  wire  axi4yank_clock; // @[UserYanker.scala 105:30]
  wire  axi4yank_reset; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_awready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_awvalid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_awid; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_in_awaddr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_awlen; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_awsize; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_awecho_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_awecho_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_wready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_wvalid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_in_wdata; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_wstrb; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_wlast; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_bready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_bvalid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_bid; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_bresp; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_becho_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_becho_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_arready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_arvalid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_arid; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_in_araddr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_arlen; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_arsize; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_arecho_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_arecho_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_rready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_rvalid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_rid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_in_rdata; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_rresp; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_recho_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_recho_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_rlast; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_awready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_awvalid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_awid; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_out_awaddr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_awlen; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_awsize; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_wready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_wvalid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_out_wdata; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_wstrb; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_wlast; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_bready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_bvalid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_bid; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_bresp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_arready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_arvalid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_arid; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_out_araddr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_arlen; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_arsize; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_rready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_rvalid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_rid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_out_rdata; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_rresp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_rlast; // @[UserYanker.scala 105:30]
  wire  axi4frag_clock; // @[Fragmenter.scala 205:30]
  wire  axi4frag_reset; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_awready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_awvalid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_awid; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_in_awaddr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_awlen; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_awsize; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_awburst; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_awecho_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_wready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_wvalid; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_in_wdata; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_wstrb; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_wlast; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_bready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_bvalid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_bid; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_bresp; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_becho_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_arready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_arvalid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_arid; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_in_araddr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_arlen; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_arsize; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_arburst; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_arecho_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_rready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_rvalid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_rid; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_in_rdata; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_rresp; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_recho_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_rlast; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_awready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_awvalid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_awid; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_out_awaddr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_awlen; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_awsize; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_awecho_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_awecho_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_wready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_wvalid; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_out_wdata; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_wstrb; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_wlast; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_bready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_bvalid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_bid; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_out_bresp; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_becho_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_becho_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_arready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_arvalid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_arid; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_out_araddr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_arlen; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_arsize; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_arecho_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_arecho_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_rready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_rvalid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_rid; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_out_rdata; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_out_rresp; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_recho_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_recho_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_rlast; // @[Fragmenter.scala 205:30]
  wire  axi4index_auto_in_awready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_awvalid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_awid; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_in_awaddr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_awlen; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_awsize; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_awburst; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_wready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_wvalid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_in_wdata; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_wstrb; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_wlast; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_bready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_bvalid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_bid; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_bresp; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_arready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_arvalid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_arid; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_in_araddr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_arlen; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_arsize; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_arburst; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_rready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_rvalid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_rid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_in_rdata; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_rresp; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_rlast; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_awready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_awvalid; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_awid; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_out_awaddr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_awlen; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_awsize; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_awburst; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_awecho_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_wready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_wvalid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_out_wdata; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_wstrb; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_wlast; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_bready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_bvalid; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_bid; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_bresp; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_becho_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_arready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_arvalid; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_arid; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_out_araddr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_arlen; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_arsize; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_arburst; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_arecho_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_rready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_rvalid; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_rid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_out_rdata; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_rresp; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_recho_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_rlast; // @[IdIndexer.scala 91:31]
  wire  axi4yank_1_clock; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_reset; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_awready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_awvalid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_in_awid; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_1_auto_in_awaddr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_1_auto_in_awlen; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_1_auto_in_awsize; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_1_auto_in_awburst; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_in_awecho_tl_state_size; // @[UserYanker.scala 105:30]
  wire [6:0] axi4yank_1_auto_in_awecho_tl_state_source; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_awecho_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_wready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_wvalid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_1_auto_in_wdata; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_1_auto_in_wstrb; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_wlast; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_bready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_bvalid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_in_bid; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_1_auto_in_bresp; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_in_becho_tl_state_size; // @[UserYanker.scala 105:30]
  wire [6:0] axi4yank_1_auto_in_becho_tl_state_source; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_becho_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_arready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_arvalid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_in_arid; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_1_auto_in_araddr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_1_auto_in_arlen; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_1_auto_in_arsize; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_1_auto_in_arburst; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_in_arecho_tl_state_size; // @[UserYanker.scala 105:30]
  wire [6:0] axi4yank_1_auto_in_arecho_tl_state_source; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_arecho_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_rready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_rvalid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_in_rid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_1_auto_in_rdata; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_1_auto_in_rresp; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_in_recho_tl_state_size; // @[UserYanker.scala 105:30]
  wire [6:0] axi4yank_1_auto_in_recho_tl_state_source; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_recho_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_in_rlast; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_awready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_awvalid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_out_awid; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_1_auto_out_awaddr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_1_auto_out_awlen; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_1_auto_out_awsize; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_1_auto_out_awburst; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_wready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_wvalid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_1_auto_out_wdata; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_1_auto_out_wstrb; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_wlast; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_bready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_bvalid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_out_bid; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_1_auto_out_bresp; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_arready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_arvalid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_out_arid; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_1_auto_out_araddr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_1_auto_out_arlen; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_1_auto_out_arsize; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_1_auto_out_arburst; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_rready; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_rvalid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_1_auto_out_rid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_1_auto_out_rdata; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_1_auto_out_rresp; // @[UserYanker.scala 105:30]
  wire  axi4yank_1_auto_out_rlast; // @[UserYanker.scala 105:30]
  wire  axi4index_1_auto_in_awready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_awvalid; // @[IdIndexer.scala 91:31]
  wire [4:0] axi4index_1_auto_in_awid; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_1_auto_in_awaddr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_1_auto_in_awlen; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_1_auto_in_awsize; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_1_auto_in_awburst; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_in_awecho_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_1_auto_in_awecho_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_wready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_wvalid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_1_auto_in_wdata; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_1_auto_in_wstrb; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_wlast; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_bready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_bvalid; // @[IdIndexer.scala 91:31]
  wire [4:0] axi4index_1_auto_in_bid; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_1_auto_in_bresp; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_in_becho_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_1_auto_in_becho_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_arready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_arvalid; // @[IdIndexer.scala 91:31]
  wire [4:0] axi4index_1_auto_in_arid; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_1_auto_in_araddr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_1_auto_in_arlen; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_1_auto_in_arsize; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_1_auto_in_arburst; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_in_arecho_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_1_auto_in_arecho_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_rready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_rvalid; // @[IdIndexer.scala 91:31]
  wire [4:0] axi4index_1_auto_in_rid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_1_auto_in_rdata; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_1_auto_in_rresp; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_in_recho_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_1_auto_in_recho_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_in_rlast; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_awready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_awvalid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_out_awid; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_1_auto_out_awaddr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_1_auto_out_awlen; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_1_auto_out_awsize; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_1_auto_out_awburst; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_out_awecho_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_1_auto_out_awecho_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_awecho_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_wready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_wvalid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_1_auto_out_wdata; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_1_auto_out_wstrb; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_wlast; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_bready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_bvalid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_out_bid; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_1_auto_out_bresp; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_out_becho_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_1_auto_out_becho_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_becho_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_arready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_arvalid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_out_arid; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_1_auto_out_araddr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_1_auto_out_arlen; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_1_auto_out_arsize; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_1_auto_out_arburst; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_out_arecho_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_1_auto_out_arecho_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_arecho_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_rready; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_rvalid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_out_rid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_1_auto_out_rdata; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_1_auto_out_rresp; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_1_auto_out_recho_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_1_auto_out_recho_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_recho_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_1_auto_out_rlast; // @[IdIndexer.scala 91:31]
  wire  tl2axi4_clock; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_reset; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_valid; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_a_bits_opcode; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_a_bits_param; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_a_bits_size; // @[ToAXI4.scala 283:29]
  wire [6:0] tl2axi4_auto_in_a_bits_source; // @[ToAXI4.scala 283:29]
  wire [31:0] tl2axi4_auto_in_a_bits_address; // @[ToAXI4.scala 283:29]
  wire [7:0] tl2axi4_auto_in_a_bits_mask; // @[ToAXI4.scala 283:29]
  wire [63:0] tl2axi4_auto_in_a_bits_data; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_bits_corrupt; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_d_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_d_valid; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_d_bits_opcode; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_d_bits_size; // @[ToAXI4.scala 283:29]
  wire [6:0] tl2axi4_auto_in_d_bits_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_d_bits_denied; // @[ToAXI4.scala 283:29]
  wire [63:0] tl2axi4_auto_in_d_bits_data; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_d_bits_corrupt; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_awready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_awvalid; // @[ToAXI4.scala 283:29]
  wire [4:0] tl2axi4_auto_out_awid; // @[ToAXI4.scala 283:29]
  wire [31:0] tl2axi4_auto_out_awaddr; // @[ToAXI4.scala 283:29]
  wire [7:0] tl2axi4_auto_out_awlen; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_out_awsize; // @[ToAXI4.scala 283:29]
  wire [1:0] tl2axi4_auto_out_awburst; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_awecho_tl_state_size; // @[ToAXI4.scala 283:29]
  wire [6:0] tl2axi4_auto_out_awecho_tl_state_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_wready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_wvalid; // @[ToAXI4.scala 283:29]
  wire [63:0] tl2axi4_auto_out_wdata; // @[ToAXI4.scala 283:29]
  wire [7:0] tl2axi4_auto_out_wstrb; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_wlast; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_bready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_bvalid; // @[ToAXI4.scala 283:29]
  wire [4:0] tl2axi4_auto_out_bid; // @[ToAXI4.scala 283:29]
  wire [1:0] tl2axi4_auto_out_bresp; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_becho_tl_state_size; // @[ToAXI4.scala 283:29]
  wire [6:0] tl2axi4_auto_out_becho_tl_state_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_arready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_arvalid; // @[ToAXI4.scala 283:29]
  wire [4:0] tl2axi4_auto_out_arid; // @[ToAXI4.scala 283:29]
  wire [31:0] tl2axi4_auto_out_araddr; // @[ToAXI4.scala 283:29]
  wire [7:0] tl2axi4_auto_out_arlen; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_out_arsize; // @[ToAXI4.scala 283:29]
  wire [1:0] tl2axi4_auto_out_arburst; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_arecho_tl_state_size; // @[ToAXI4.scala 283:29]
  wire [6:0] tl2axi4_auto_out_arecho_tl_state_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_rready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_rvalid; // @[ToAXI4.scala 283:29]
  wire [4:0] tl2axi4_auto_out_rid; // @[ToAXI4.scala 283:29]
  wire [63:0] tl2axi4_auto_out_rdata; // @[ToAXI4.scala 283:29]
  wire [1:0] tl2axi4_auto_out_rresp; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_recho_tl_state_size; // @[ToAXI4.scala 283:29]
  wire [6:0] tl2axi4_auto_out_recho_tl_state_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_rlast; // @[ToAXI4.scala 283:29]
  wire  err_clock; // @[ChipLinkBridge.scala 150:23]
  wire  err_reset; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_a_ready; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_a_valid; // @[ChipLinkBridge.scala 150:23]
  wire [2:0] err_auto_in_a_bits_opcode; // @[ChipLinkBridge.scala 150:23]
  wire [2:0] err_auto_in_a_bits_param; // @[ChipLinkBridge.scala 150:23]
  wire [2:0] err_auto_in_a_bits_size; // @[ChipLinkBridge.scala 150:23]
  wire [6:0] err_auto_in_a_bits_source; // @[ChipLinkBridge.scala 150:23]
  wire [12:0] err_auto_in_a_bits_address; // @[ChipLinkBridge.scala 150:23]
  wire [3:0] err_auto_in_a_bits_mask; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_a_bits_corrupt; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_c_ready; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_c_valid; // @[ChipLinkBridge.scala 150:23]
  wire [2:0] err_auto_in_c_bits_opcode; // @[ChipLinkBridge.scala 150:23]
  wire [2:0] err_auto_in_c_bits_param; // @[ChipLinkBridge.scala 150:23]
  wire [2:0] err_auto_in_c_bits_size; // @[ChipLinkBridge.scala 150:23]
  wire [6:0] err_auto_in_c_bits_source; // @[ChipLinkBridge.scala 150:23]
  wire [12:0] err_auto_in_c_bits_address; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_d_ready; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_d_valid; // @[ChipLinkBridge.scala 150:23]
  wire [2:0] err_auto_in_d_bits_opcode; // @[ChipLinkBridge.scala 150:23]
  wire [1:0] err_auto_in_d_bits_param; // @[ChipLinkBridge.scala 150:23]
  wire [2:0] err_auto_in_d_bits_size; // @[ChipLinkBridge.scala 150:23]
  wire [6:0] err_auto_in_d_bits_source; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_d_bits_denied; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_d_bits_corrupt; // @[ChipLinkBridge.scala 150:23]
  wire  err_auto_in_e_valid; // @[ChipLinkBridge.scala 150:23]
  wire  atomics_clock; // @[AtomicAutomata.scala 283:29]
  wire  atomics_reset; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_a_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_a_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_a_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_a_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_a_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_in_a_bits_source; // @[AtomicAutomata.scala 283:29]
  wire [31:0] atomics_auto_in_a_bits_address; // @[AtomicAutomata.scala 283:29]
  wire [7:0] atomics_auto_in_a_bits_mask; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_in_a_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_c_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_c_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_c_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_c_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_c_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_in_c_bits_source; // @[AtomicAutomata.scala 283:29]
  wire [31:0] atomics_auto_in_c_bits_address; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_d_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [1:0] atomics_auto_in_d_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_d_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_in_d_bits_source; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_bits_denied; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_in_d_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_bits_corrupt; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_e_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_e_valid; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_e_bits_sink; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_a_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_a_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_a_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_a_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_a_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_out_a_bits_source; // @[AtomicAutomata.scala 283:29]
  wire [31:0] atomics_auto_out_a_bits_address; // @[AtomicAutomata.scala 283:29]
  wire [7:0] atomics_auto_out_a_bits_mask; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_out_a_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_a_bits_corrupt; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_c_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_c_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_c_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_c_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_c_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_out_c_bits_source; // @[AtomicAutomata.scala 283:29]
  wire [31:0] atomics_auto_out_c_bits_address; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_d_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [1:0] atomics_auto_out_d_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_d_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_out_d_bits_source; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_bits_denied; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_out_d_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_bits_corrupt; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_e_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_e_valid; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_e_bits_sink; // @[AtomicAutomata.scala 283:29]
  wire  fixer_1_clock; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_reset; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_in_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_in_a_bits_param; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_in_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [6:0] fixer_1_auto_in_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_1_auto_in_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_1_auto_in_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_1_auto_in_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_c_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_c_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_in_c_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_in_c_bits_param; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_in_c_bits_size; // @[FIFOFixer.scala 144:27]
  wire [6:0] fixer_1_auto_in_c_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_1_auto_in_c_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_in_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [1:0] fixer_1_auto_in_d_bits_param; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_in_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [6:0] fixer_1_auto_in_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_1_auto_in_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_e_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_e_valid; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_in_e_bits_sink; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_out_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_out_a_bits_param; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_out_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [6:0] fixer_1_auto_out_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_1_auto_out_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_1_auto_out_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_1_auto_out_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_c_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_c_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_out_c_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_out_c_bits_param; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_out_c_bits_size; // @[FIFOFixer.scala 144:27]
  wire [6:0] fixer_1_auto_out_c_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_1_auto_out_c_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_out_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [1:0] fixer_1_auto_out_d_bits_param; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_1_auto_out_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [6:0] fixer_1_auto_out_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_1_auto_out_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_e_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_e_valid; // @[FIFOFixer.scala 144:27]
  wire  fixer_1_auto_out_e_bits_sink; // @[FIFOFixer.scala 144:27]
  wire  hints_clock; // @[HintHandler.scala 119:27]
  wire  hints_reset; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_a_ready; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_a_valid; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_in_a_bits_opcode; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_in_a_bits_param; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_in_a_bits_size; // @[HintHandler.scala 119:27]
  wire [5:0] hints_auto_in_a_bits_source; // @[HintHandler.scala 119:27]
  wire [31:0] hints_auto_in_a_bits_address; // @[HintHandler.scala 119:27]
  wire [7:0] hints_auto_in_a_bits_mask; // @[HintHandler.scala 119:27]
  wire [63:0] hints_auto_in_a_bits_data; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_c_ready; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_c_valid; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_in_c_bits_opcode; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_in_c_bits_param; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_in_c_bits_size; // @[HintHandler.scala 119:27]
  wire [5:0] hints_auto_in_c_bits_source; // @[HintHandler.scala 119:27]
  wire [31:0] hints_auto_in_c_bits_address; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_d_ready; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_d_valid; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_in_d_bits_opcode; // @[HintHandler.scala 119:27]
  wire [1:0] hints_auto_in_d_bits_param; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_in_d_bits_size; // @[HintHandler.scala 119:27]
  wire [5:0] hints_auto_in_d_bits_source; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_d_bits_denied; // @[HintHandler.scala 119:27]
  wire [63:0] hints_auto_in_d_bits_data; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_d_bits_corrupt; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_e_ready; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_e_valid; // @[HintHandler.scala 119:27]
  wire  hints_auto_in_e_bits_sink; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_a_ready; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_a_valid; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_out_a_bits_opcode; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_out_a_bits_param; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_out_a_bits_size; // @[HintHandler.scala 119:27]
  wire [6:0] hints_auto_out_a_bits_source; // @[HintHandler.scala 119:27]
  wire [31:0] hints_auto_out_a_bits_address; // @[HintHandler.scala 119:27]
  wire [7:0] hints_auto_out_a_bits_mask; // @[HintHandler.scala 119:27]
  wire [63:0] hints_auto_out_a_bits_data; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_c_ready; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_c_valid; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_out_c_bits_opcode; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_out_c_bits_param; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_out_c_bits_size; // @[HintHandler.scala 119:27]
  wire [6:0] hints_auto_out_c_bits_source; // @[HintHandler.scala 119:27]
  wire [31:0] hints_auto_out_c_bits_address; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_d_ready; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_d_valid; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_out_d_bits_opcode; // @[HintHandler.scala 119:27]
  wire [1:0] hints_auto_out_d_bits_param; // @[HintHandler.scala 119:27]
  wire [2:0] hints_auto_out_d_bits_size; // @[HintHandler.scala 119:27]
  wire [6:0] hints_auto_out_d_bits_source; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_d_bits_denied; // @[HintHandler.scala 119:27]
  wire [63:0] hints_auto_out_d_bits_data; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_d_bits_corrupt; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_e_ready; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_e_valid; // @[HintHandler.scala 119:27]
  wire  hints_auto_out_e_bits_sink; // @[HintHandler.scala 119:27]
  wire  widget_1_clock; // @[WidthWidget.scala 219:28]
  wire  widget_1_reset; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_a_ready; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_a_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_in_a_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_in_a_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_in_a_bits_size; // @[WidthWidget.scala 219:28]
  wire [5:0] widget_1_auto_in_a_bits_source; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_1_auto_in_a_bits_address; // @[WidthWidget.scala 219:28]
  wire [3:0] widget_1_auto_in_a_bits_mask; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_1_auto_in_a_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_c_ready; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_c_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_in_c_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_in_c_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_in_c_bits_size; // @[WidthWidget.scala 219:28]
  wire [5:0] widget_1_auto_in_c_bits_source; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_1_auto_in_c_bits_address; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_d_ready; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_d_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_in_d_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [1:0] widget_1_auto_in_d_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_in_d_bits_size; // @[WidthWidget.scala 219:28]
  wire [5:0] widget_1_auto_in_d_bits_source; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_d_bits_denied; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_1_auto_in_d_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_d_bits_corrupt; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_e_ready; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_e_valid; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_in_e_bits_sink; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_a_ready; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_a_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_out_a_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_out_a_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_out_a_bits_size; // @[WidthWidget.scala 219:28]
  wire [5:0] widget_1_auto_out_a_bits_source; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_1_auto_out_a_bits_address; // @[WidthWidget.scala 219:28]
  wire [7:0] widget_1_auto_out_a_bits_mask; // @[WidthWidget.scala 219:28]
  wire [63:0] widget_1_auto_out_a_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_c_ready; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_c_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_out_c_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_out_c_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_out_c_bits_size; // @[WidthWidget.scala 219:28]
  wire [5:0] widget_1_auto_out_c_bits_source; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_1_auto_out_c_bits_address; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_d_ready; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_d_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_out_d_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [1:0] widget_1_auto_out_d_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_1_auto_out_d_bits_size; // @[WidthWidget.scala 219:28]
  wire [5:0] widget_1_auto_out_d_bits_source; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_d_bits_denied; // @[WidthWidget.scala 219:28]
  wire [63:0] widget_1_auto_out_d_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_d_bits_corrupt; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_e_ready; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_e_valid; // @[WidthWidget.scala 219:28]
  wire  widget_1_auto_out_e_bits_sink; // @[WidthWidget.scala 219:28]
  wire  widget_2_clock; // @[WidthWidget.scala 219:28]
  wire  widget_2_reset; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_a_ready; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_a_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_in_a_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_in_a_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_in_a_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_2_auto_in_a_bits_source; // @[WidthWidget.scala 219:28]
  wire [12:0] widget_2_auto_in_a_bits_address; // @[WidthWidget.scala 219:28]
  wire [7:0] widget_2_auto_in_a_bits_mask; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_a_bits_corrupt; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_c_ready; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_c_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_in_c_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_in_c_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_in_c_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_2_auto_in_c_bits_source; // @[WidthWidget.scala 219:28]
  wire [12:0] widget_2_auto_in_c_bits_address; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_d_ready; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_d_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_in_d_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [1:0] widget_2_auto_in_d_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_in_d_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_2_auto_in_d_bits_source; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_d_bits_denied; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_d_bits_corrupt; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_in_e_valid; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_a_ready; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_a_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_out_a_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_out_a_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_out_a_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_2_auto_out_a_bits_source; // @[WidthWidget.scala 219:28]
  wire [12:0] widget_2_auto_out_a_bits_address; // @[WidthWidget.scala 219:28]
  wire [3:0] widget_2_auto_out_a_bits_mask; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_a_bits_corrupt; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_c_ready; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_c_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_out_c_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_out_c_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_out_c_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_2_auto_out_c_bits_source; // @[WidthWidget.scala 219:28]
  wire [12:0] widget_2_auto_out_c_bits_address; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_d_ready; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_d_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_out_d_bits_opcode; // @[WidthWidget.scala 219:28]
  wire [1:0] widget_2_auto_out_d_bits_param; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_2_auto_out_d_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_2_auto_out_d_bits_source; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_d_bits_denied; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_d_bits_corrupt; // @[WidthWidget.scala 219:28]
  wire  widget_2_auto_out_e_valid; // @[WidthWidget.scala 219:28]
  TLXbar xbar ( // @[Xbar.scala 142:26]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .auto_in_a_ready(xbar_auto_in_a_ready),
    .auto_in_a_valid(xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(xbar_auto_in_a_bits_corrupt),
    .auto_in_c_ready(xbar_auto_in_c_ready),
    .auto_in_c_valid(xbar_auto_in_c_valid),
    .auto_in_c_bits_opcode(xbar_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(xbar_auto_in_c_bits_param),
    .auto_in_c_bits_size(xbar_auto_in_c_bits_size),
    .auto_in_c_bits_source(xbar_auto_in_c_bits_source),
    .auto_in_c_bits_address(xbar_auto_in_c_bits_address),
    .auto_in_d_ready(xbar_auto_in_d_ready),
    .auto_in_d_valid(xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_auto_in_d_bits_source),
    .auto_in_d_bits_denied(xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_auto_in_d_bits_corrupt),
    .auto_in_e_ready(xbar_auto_in_e_ready),
    .auto_in_e_valid(xbar_auto_in_e_valid),
    .auto_in_e_bits_sink(xbar_auto_in_e_bits_sink),
    .auto_out_1_a_ready(xbar_auto_out_1_a_ready),
    .auto_out_1_a_valid(xbar_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(xbar_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_param(xbar_auto_out_1_a_bits_param),
    .auto_out_1_a_bits_size(xbar_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(xbar_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(xbar_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_mask(xbar_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_corrupt(xbar_auto_out_1_a_bits_corrupt),
    .auto_out_1_c_ready(xbar_auto_out_1_c_ready),
    .auto_out_1_c_valid(xbar_auto_out_1_c_valid),
    .auto_out_1_c_bits_opcode(xbar_auto_out_1_c_bits_opcode),
    .auto_out_1_c_bits_param(xbar_auto_out_1_c_bits_param),
    .auto_out_1_c_bits_size(xbar_auto_out_1_c_bits_size),
    .auto_out_1_c_bits_source(xbar_auto_out_1_c_bits_source),
    .auto_out_1_c_bits_address(xbar_auto_out_1_c_bits_address),
    .auto_out_1_d_ready(xbar_auto_out_1_d_ready),
    .auto_out_1_d_valid(xbar_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(xbar_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_param(xbar_auto_out_1_d_bits_param),
    .auto_out_1_d_bits_size(xbar_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(xbar_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_denied(xbar_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_corrupt(xbar_auto_out_1_d_bits_corrupt),
    .auto_out_1_e_valid(xbar_auto_out_1_e_valid),
    .auto_out_0_a_ready(xbar_auto_out_0_a_ready),
    .auto_out_0_a_valid(xbar_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(xbar_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_param(xbar_auto_out_0_a_bits_param),
    .auto_out_0_a_bits_size(xbar_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(xbar_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(xbar_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_mask(xbar_auto_out_0_a_bits_mask),
    .auto_out_0_a_bits_data(xbar_auto_out_0_a_bits_data),
    .auto_out_0_a_bits_corrupt(xbar_auto_out_0_a_bits_corrupt),
    .auto_out_0_d_ready(xbar_auto_out_0_d_ready),
    .auto_out_0_d_valid(xbar_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(xbar_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_size(xbar_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(xbar_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_denied(xbar_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(xbar_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(xbar_auto_out_0_d_bits_corrupt)
  );
  TLXbar_1 xbar_1 ( // @[Xbar.scala 142:26]
    .clock(xbar_1_clock),
    .reset(xbar_1_reset),
    .auto_in_a_ready(xbar_1_auto_in_a_ready),
    .auto_in_a_valid(xbar_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(xbar_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_1_auto_in_a_bits_data),
    .auto_in_d_ready(xbar_1_auto_in_d_ready),
    .auto_in_d_valid(xbar_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_1_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_1_auto_in_d_bits_source),
    .auto_in_d_bits_sink(xbar_1_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(xbar_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_1_auto_in_d_bits_corrupt),
    .auto_out_1_a_ready(xbar_1_auto_out_1_a_ready),
    .auto_out_1_a_valid(xbar_1_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(xbar_1_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_size(xbar_1_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(xbar_1_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(xbar_1_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_mask(xbar_1_auto_out_1_a_bits_mask),
    .auto_out_1_d_ready(xbar_1_auto_out_1_d_ready),
    .auto_out_1_d_valid(xbar_1_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(xbar_1_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_size(xbar_1_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(xbar_1_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_denied(xbar_1_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_corrupt(xbar_1_auto_out_1_d_bits_corrupt),
    .auto_out_0_a_ready(xbar_1_auto_out_0_a_ready),
    .auto_out_0_a_valid(xbar_1_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(xbar_1_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_size(xbar_1_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(xbar_1_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(xbar_1_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_mask(xbar_1_auto_out_0_a_bits_mask),
    .auto_out_0_a_bits_data(xbar_1_auto_out_0_a_bits_data),
    .auto_out_0_d_ready(xbar_1_auto_out_0_d_ready),
    .auto_out_0_d_valid(xbar_1_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(xbar_1_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_param(xbar_1_auto_out_0_d_bits_param),
    .auto_out_0_d_bits_size(xbar_1_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(xbar_1_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_sink(xbar_1_auto_out_0_d_bits_sink),
    .auto_out_0_d_bits_denied(xbar_1_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(xbar_1_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(xbar_1_auto_out_0_d_bits_corrupt)
  );
  TLError ferr ( // @[ChipLinkBridge.scala 31:24]
    .clock(ferr_clock),
    .reset(ferr_reset),
    .auto_in_a_ready(ferr_auto_in_a_ready),
    .auto_in_a_valid(ferr_auto_in_a_valid),
    .auto_in_a_bits_opcode(ferr_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(ferr_auto_in_a_bits_size),
    .auto_in_a_bits_source(ferr_auto_in_a_bits_source),
    .auto_in_a_bits_address(ferr_auto_in_a_bits_address),
    .auto_in_a_bits_mask(ferr_auto_in_a_bits_mask),
    .auto_in_d_ready(ferr_auto_in_d_ready),
    .auto_in_d_valid(ferr_auto_in_d_valid),
    .auto_in_d_bits_opcode(ferr_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(ferr_auto_in_d_bits_size),
    .auto_in_d_bits_source(ferr_auto_in_d_bits_source),
    .auto_in_d_bits_denied(ferr_auto_in_d_bits_denied),
    .auto_in_d_bits_corrupt(ferr_auto_in_d_bits_corrupt)
  );
  ChipLink chiplink ( // @[ChipLinkBridge.scala 39:28]
    .clock(chiplink_clock),
    .reset(chiplink_reset),
    .auto_mbypass_out_a_ready(chiplink_auto_mbypass_out_a_ready),
    .auto_mbypass_out_a_valid(chiplink_auto_mbypass_out_a_valid),
    .auto_mbypass_out_a_bits_opcode(chiplink_auto_mbypass_out_a_bits_opcode),
    .auto_mbypass_out_a_bits_param(chiplink_auto_mbypass_out_a_bits_param),
    .auto_mbypass_out_a_bits_size(chiplink_auto_mbypass_out_a_bits_size),
    .auto_mbypass_out_a_bits_source(chiplink_auto_mbypass_out_a_bits_source),
    .auto_mbypass_out_a_bits_address(chiplink_auto_mbypass_out_a_bits_address),
    .auto_mbypass_out_a_bits_mask(chiplink_auto_mbypass_out_a_bits_mask),
    .auto_mbypass_out_a_bits_data(chiplink_auto_mbypass_out_a_bits_data),
    .auto_mbypass_out_c_ready(chiplink_auto_mbypass_out_c_ready),
    .auto_mbypass_out_c_valid(chiplink_auto_mbypass_out_c_valid),
    .auto_mbypass_out_c_bits_opcode(chiplink_auto_mbypass_out_c_bits_opcode),
    .auto_mbypass_out_c_bits_param(chiplink_auto_mbypass_out_c_bits_param),
    .auto_mbypass_out_c_bits_size(chiplink_auto_mbypass_out_c_bits_size),
    .auto_mbypass_out_c_bits_source(chiplink_auto_mbypass_out_c_bits_source),
    .auto_mbypass_out_c_bits_address(chiplink_auto_mbypass_out_c_bits_address),
    .auto_mbypass_out_d_ready(chiplink_auto_mbypass_out_d_ready),
    .auto_mbypass_out_d_valid(chiplink_auto_mbypass_out_d_valid),
    .auto_mbypass_out_d_bits_opcode(chiplink_auto_mbypass_out_d_bits_opcode),
    .auto_mbypass_out_d_bits_param(chiplink_auto_mbypass_out_d_bits_param),
    .auto_mbypass_out_d_bits_size(chiplink_auto_mbypass_out_d_bits_size),
    .auto_mbypass_out_d_bits_source(chiplink_auto_mbypass_out_d_bits_source),
    .auto_mbypass_out_d_bits_denied(chiplink_auto_mbypass_out_d_bits_denied),
    .auto_mbypass_out_d_bits_data(chiplink_auto_mbypass_out_d_bits_data),
    .auto_mbypass_out_d_bits_corrupt(chiplink_auto_mbypass_out_d_bits_corrupt),
    .auto_mbypass_out_e_ready(chiplink_auto_mbypass_out_e_ready),
    .auto_mbypass_out_e_valid(chiplink_auto_mbypass_out_e_valid),
    .auto_mbypass_out_e_bits_sink(chiplink_auto_mbypass_out_e_bits_sink),
    .auto_sbypass_node_in_in_a_ready(chiplink_auto_sbypass_node_in_in_a_ready),
    .auto_sbypass_node_in_in_a_valid(chiplink_auto_sbypass_node_in_in_a_valid),
    .auto_sbypass_node_in_in_a_bits_opcode(chiplink_auto_sbypass_node_in_in_a_bits_opcode),
    .auto_sbypass_node_in_in_a_bits_size(chiplink_auto_sbypass_node_in_in_a_bits_size),
    .auto_sbypass_node_in_in_a_bits_source(chiplink_auto_sbypass_node_in_in_a_bits_source),
    .auto_sbypass_node_in_in_a_bits_address(chiplink_auto_sbypass_node_in_in_a_bits_address),
    .auto_sbypass_node_in_in_a_bits_mask(chiplink_auto_sbypass_node_in_in_a_bits_mask),
    .auto_sbypass_node_in_in_a_bits_data(chiplink_auto_sbypass_node_in_in_a_bits_data),
    .auto_sbypass_node_in_in_d_ready(chiplink_auto_sbypass_node_in_in_d_ready),
    .auto_sbypass_node_in_in_d_valid(chiplink_auto_sbypass_node_in_in_d_valid),
    .auto_sbypass_node_in_in_d_bits_opcode(chiplink_auto_sbypass_node_in_in_d_bits_opcode),
    .auto_sbypass_node_in_in_d_bits_param(chiplink_auto_sbypass_node_in_in_d_bits_param),
    .auto_sbypass_node_in_in_d_bits_size(chiplink_auto_sbypass_node_in_in_d_bits_size),
    .auto_sbypass_node_in_in_d_bits_source(chiplink_auto_sbypass_node_in_in_d_bits_source),
    .auto_sbypass_node_in_in_d_bits_sink(chiplink_auto_sbypass_node_in_in_d_bits_sink),
    .auto_sbypass_node_in_in_d_bits_denied(chiplink_auto_sbypass_node_in_in_d_bits_denied),
    .auto_sbypass_node_in_in_d_bits_data(chiplink_auto_sbypass_node_in_in_d_bits_data),
    .auto_sbypass_node_in_in_d_bits_corrupt(chiplink_auto_sbypass_node_in_in_d_bits_corrupt),
    .auto_io_out_c2b_clk(chiplink_auto_io_out_c2b_clk),
    .auto_io_out_c2b_rst(chiplink_auto_io_out_c2b_rst),
    .auto_io_out_c2b_send(chiplink_auto_io_out_c2b_send),
    .auto_io_out_c2b_data(chiplink_auto_io_out_c2b_data),
    .auto_io_out_b2c_clk(chiplink_auto_io_out_b2c_clk),
    .auto_io_out_b2c_rst(chiplink_auto_io_out_b2c_rst),
    .auto_io_out_b2c_send(chiplink_auto_io_out_b2c_send),
    .auto_io_out_b2c_data(chiplink_auto_io_out_b2c_data)
  );
  TLFIFOFixer fixer ( // @[FIFOFixer.scala 144:27]
    .clock(fixer_clock),
    .reset(fixer_reset),
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fixer_auto_in_d_bits_param),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fixer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fixer_auto_out_d_bits_param),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fixer_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt)
  );
  TLWidthWidget widget ( // @[WidthWidget.scala 219:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_auto_in_a_bits_data),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(widget_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_auto_in_d_bits_source),
    .auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_auto_out_a_bits_data),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
  );
  AXI4ToTL axi42tl ( // @[ToTL.scala 216:29]
    .clock(axi42tl_clock),
    .reset(axi42tl_reset),
    .auto_in_awready(axi42tl_auto_in_awready),
    .auto_in_awvalid(axi42tl_auto_in_awvalid),
    .auto_in_awid(axi42tl_auto_in_awid),
    .auto_in_awaddr(axi42tl_auto_in_awaddr),
    .auto_in_awlen(axi42tl_auto_in_awlen),
    .auto_in_awsize(axi42tl_auto_in_awsize),
    .auto_in_wready(axi42tl_auto_in_wready),
    .auto_in_wvalid(axi42tl_auto_in_wvalid),
    .auto_in_wdata(axi42tl_auto_in_wdata),
    .auto_in_wstrb(axi42tl_auto_in_wstrb),
    .auto_in_wlast(axi42tl_auto_in_wlast),
    .auto_in_bready(axi42tl_auto_in_bready),
    .auto_in_bvalid(axi42tl_auto_in_bvalid),
    .auto_in_bid(axi42tl_auto_in_bid),
    .auto_in_bresp(axi42tl_auto_in_bresp),
    .auto_in_arready(axi42tl_auto_in_arready),
    .auto_in_arvalid(axi42tl_auto_in_arvalid),
    .auto_in_arid(axi42tl_auto_in_arid),
    .auto_in_araddr(axi42tl_auto_in_araddr),
    .auto_in_arlen(axi42tl_auto_in_arlen),
    .auto_in_arsize(axi42tl_auto_in_arsize),
    .auto_in_rready(axi42tl_auto_in_rready),
    .auto_in_rvalid(axi42tl_auto_in_rvalid),
    .auto_in_rid(axi42tl_auto_in_rid),
    .auto_in_rdata(axi42tl_auto_in_rdata),
    .auto_in_rresp(axi42tl_auto_in_rresp),
    .auto_in_rlast(axi42tl_auto_in_rlast),
    .auto_out_a_ready(axi42tl_auto_out_a_ready),
    .auto_out_a_valid(axi42tl_auto_out_a_valid),
    .auto_out_a_bits_opcode(axi42tl_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(axi42tl_auto_out_a_bits_size),
    .auto_out_a_bits_source(axi42tl_auto_out_a_bits_source),
    .auto_out_a_bits_address(axi42tl_auto_out_a_bits_address),
    .auto_out_a_bits_mask(axi42tl_auto_out_a_bits_mask),
    .auto_out_a_bits_data(axi42tl_auto_out_a_bits_data),
    .auto_out_d_ready(axi42tl_auto_out_d_ready),
    .auto_out_d_valid(axi42tl_auto_out_d_valid),
    .auto_out_d_bits_opcode(axi42tl_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(axi42tl_auto_out_d_bits_size),
    .auto_out_d_bits_source(axi42tl_auto_out_d_bits_source),
    .auto_out_d_bits_denied(axi42tl_auto_out_d_bits_denied),
    .auto_out_d_bits_data(axi42tl_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(axi42tl_auto_out_d_bits_corrupt)
  );
  AXI4UserYanker axi4yank ( // @[UserYanker.scala 105:30]
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_awready(axi4yank_auto_in_awready),
    .auto_in_awvalid(axi4yank_auto_in_awvalid),
    .auto_in_awid(axi4yank_auto_in_awid),
    .auto_in_awaddr(axi4yank_auto_in_awaddr),
    .auto_in_awlen(axi4yank_auto_in_awlen),
    .auto_in_awsize(axi4yank_auto_in_awsize),
    .auto_in_awecho_extra_id(axi4yank_auto_in_awecho_extra_id),
    .auto_in_awecho_real_last(axi4yank_auto_in_awecho_real_last),
    .auto_in_wready(axi4yank_auto_in_wready),
    .auto_in_wvalid(axi4yank_auto_in_wvalid),
    .auto_in_wdata(axi4yank_auto_in_wdata),
    .auto_in_wstrb(axi4yank_auto_in_wstrb),
    .auto_in_wlast(axi4yank_auto_in_wlast),
    .auto_in_bready(axi4yank_auto_in_bready),
    .auto_in_bvalid(axi4yank_auto_in_bvalid),
    .auto_in_bid(axi4yank_auto_in_bid),
    .auto_in_bresp(axi4yank_auto_in_bresp),
    .auto_in_becho_extra_id(axi4yank_auto_in_becho_extra_id),
    .auto_in_becho_real_last(axi4yank_auto_in_becho_real_last),
    .auto_in_arready(axi4yank_auto_in_arready),
    .auto_in_arvalid(axi4yank_auto_in_arvalid),
    .auto_in_arid(axi4yank_auto_in_arid),
    .auto_in_araddr(axi4yank_auto_in_araddr),
    .auto_in_arlen(axi4yank_auto_in_arlen),
    .auto_in_arsize(axi4yank_auto_in_arsize),
    .auto_in_arecho_extra_id(axi4yank_auto_in_arecho_extra_id),
    .auto_in_arecho_real_last(axi4yank_auto_in_arecho_real_last),
    .auto_in_rready(axi4yank_auto_in_rready),
    .auto_in_rvalid(axi4yank_auto_in_rvalid),
    .auto_in_rid(axi4yank_auto_in_rid),
    .auto_in_rdata(axi4yank_auto_in_rdata),
    .auto_in_rresp(axi4yank_auto_in_rresp),
    .auto_in_recho_extra_id(axi4yank_auto_in_recho_extra_id),
    .auto_in_recho_real_last(axi4yank_auto_in_recho_real_last),
    .auto_in_rlast(axi4yank_auto_in_rlast),
    .auto_out_awready(axi4yank_auto_out_awready),
    .auto_out_awvalid(axi4yank_auto_out_awvalid),
    .auto_out_awid(axi4yank_auto_out_awid),
    .auto_out_awaddr(axi4yank_auto_out_awaddr),
    .auto_out_awlen(axi4yank_auto_out_awlen),
    .auto_out_awsize(axi4yank_auto_out_awsize),
    .auto_out_wready(axi4yank_auto_out_wready),
    .auto_out_wvalid(axi4yank_auto_out_wvalid),
    .auto_out_wdata(axi4yank_auto_out_wdata),
    .auto_out_wstrb(axi4yank_auto_out_wstrb),
    .auto_out_wlast(axi4yank_auto_out_wlast),
    .auto_out_bready(axi4yank_auto_out_bready),
    .auto_out_bvalid(axi4yank_auto_out_bvalid),
    .auto_out_bid(axi4yank_auto_out_bid),
    .auto_out_bresp(axi4yank_auto_out_bresp),
    .auto_out_arready(axi4yank_auto_out_arready),
    .auto_out_arvalid(axi4yank_auto_out_arvalid),
    .auto_out_arid(axi4yank_auto_out_arid),
    .auto_out_araddr(axi4yank_auto_out_araddr),
    .auto_out_arlen(axi4yank_auto_out_arlen),
    .auto_out_arsize(axi4yank_auto_out_arsize),
    .auto_out_rready(axi4yank_auto_out_rready),
    .auto_out_rvalid(axi4yank_auto_out_rvalid),
    .auto_out_rid(axi4yank_auto_out_rid),
    .auto_out_rdata(axi4yank_auto_out_rdata),
    .auto_out_rresp(axi4yank_auto_out_rresp),
    .auto_out_rlast(axi4yank_auto_out_rlast)
  );
  AXI4Fragmenter axi4frag ( // @[Fragmenter.scala 205:30]
    .clock(axi4frag_clock),
    .reset(axi4frag_reset),
    .auto_in_awready(axi4frag_auto_in_awready),
    .auto_in_awvalid(axi4frag_auto_in_awvalid),
    .auto_in_awid(axi4frag_auto_in_awid),
    .auto_in_awaddr(axi4frag_auto_in_awaddr),
    .auto_in_awlen(axi4frag_auto_in_awlen),
    .auto_in_awsize(axi4frag_auto_in_awsize),
    .auto_in_awburst(axi4frag_auto_in_awburst),
    .auto_in_awecho_extra_id(axi4frag_auto_in_awecho_extra_id),
    .auto_in_wready(axi4frag_auto_in_wready),
    .auto_in_wvalid(axi4frag_auto_in_wvalid),
    .auto_in_wdata(axi4frag_auto_in_wdata),
    .auto_in_wstrb(axi4frag_auto_in_wstrb),
    .auto_in_wlast(axi4frag_auto_in_wlast),
    .auto_in_bready(axi4frag_auto_in_bready),
    .auto_in_bvalid(axi4frag_auto_in_bvalid),
    .auto_in_bid(axi4frag_auto_in_bid),
    .auto_in_bresp(axi4frag_auto_in_bresp),
    .auto_in_becho_extra_id(axi4frag_auto_in_becho_extra_id),
    .auto_in_arready(axi4frag_auto_in_arready),
    .auto_in_arvalid(axi4frag_auto_in_arvalid),
    .auto_in_arid(axi4frag_auto_in_arid),
    .auto_in_araddr(axi4frag_auto_in_araddr),
    .auto_in_arlen(axi4frag_auto_in_arlen),
    .auto_in_arsize(axi4frag_auto_in_arsize),
    .auto_in_arburst(axi4frag_auto_in_arburst),
    .auto_in_arecho_extra_id(axi4frag_auto_in_arecho_extra_id),
    .auto_in_rready(axi4frag_auto_in_rready),
    .auto_in_rvalid(axi4frag_auto_in_rvalid),
    .auto_in_rid(axi4frag_auto_in_rid),
    .auto_in_rdata(axi4frag_auto_in_rdata),
    .auto_in_rresp(axi4frag_auto_in_rresp),
    .auto_in_recho_extra_id(axi4frag_auto_in_recho_extra_id),
    .auto_in_rlast(axi4frag_auto_in_rlast),
    .auto_out_awready(axi4frag_auto_out_awready),
    .auto_out_awvalid(axi4frag_auto_out_awvalid),
    .auto_out_awid(axi4frag_auto_out_awid),
    .auto_out_awaddr(axi4frag_auto_out_awaddr),
    .auto_out_awlen(axi4frag_auto_out_awlen),
    .auto_out_awsize(axi4frag_auto_out_awsize),
    .auto_out_awecho_extra_id(axi4frag_auto_out_awecho_extra_id),
    .auto_out_awecho_real_last(axi4frag_auto_out_awecho_real_last),
    .auto_out_wready(axi4frag_auto_out_wready),
    .auto_out_wvalid(axi4frag_auto_out_wvalid),
    .auto_out_wdata(axi4frag_auto_out_wdata),
    .auto_out_wstrb(axi4frag_auto_out_wstrb),
    .auto_out_wlast(axi4frag_auto_out_wlast),
    .auto_out_bready(axi4frag_auto_out_bready),
    .auto_out_bvalid(axi4frag_auto_out_bvalid),
    .auto_out_bid(axi4frag_auto_out_bid),
    .auto_out_bresp(axi4frag_auto_out_bresp),
    .auto_out_becho_extra_id(axi4frag_auto_out_becho_extra_id),
    .auto_out_becho_real_last(axi4frag_auto_out_becho_real_last),
    .auto_out_arready(axi4frag_auto_out_arready),
    .auto_out_arvalid(axi4frag_auto_out_arvalid),
    .auto_out_arid(axi4frag_auto_out_arid),
    .auto_out_araddr(axi4frag_auto_out_araddr),
    .auto_out_arlen(axi4frag_auto_out_arlen),
    .auto_out_arsize(axi4frag_auto_out_arsize),
    .auto_out_arecho_extra_id(axi4frag_auto_out_arecho_extra_id),
    .auto_out_arecho_real_last(axi4frag_auto_out_arecho_real_last),
    .auto_out_rready(axi4frag_auto_out_rready),
    .auto_out_rvalid(axi4frag_auto_out_rvalid),
    .auto_out_rid(axi4frag_auto_out_rid),
    .auto_out_rdata(axi4frag_auto_out_rdata),
    .auto_out_rresp(axi4frag_auto_out_rresp),
    .auto_out_recho_extra_id(axi4frag_auto_out_recho_extra_id),
    .auto_out_recho_real_last(axi4frag_auto_out_recho_real_last),
    .auto_out_rlast(axi4frag_auto_out_rlast)
  );
  AXI4IdIndexer axi4index ( // @[IdIndexer.scala 91:31]
    .auto_in_awready(axi4index_auto_in_awready),
    .auto_in_awvalid(axi4index_auto_in_awvalid),
    .auto_in_awid(axi4index_auto_in_awid),
    .auto_in_awaddr(axi4index_auto_in_awaddr),
    .auto_in_awlen(axi4index_auto_in_awlen),
    .auto_in_awsize(axi4index_auto_in_awsize),
    .auto_in_awburst(axi4index_auto_in_awburst),
    .auto_in_wready(axi4index_auto_in_wready),
    .auto_in_wvalid(axi4index_auto_in_wvalid),
    .auto_in_wdata(axi4index_auto_in_wdata),
    .auto_in_wstrb(axi4index_auto_in_wstrb),
    .auto_in_wlast(axi4index_auto_in_wlast),
    .auto_in_bready(axi4index_auto_in_bready),
    .auto_in_bvalid(axi4index_auto_in_bvalid),
    .auto_in_bid(axi4index_auto_in_bid),
    .auto_in_bresp(axi4index_auto_in_bresp),
    .auto_in_arready(axi4index_auto_in_arready),
    .auto_in_arvalid(axi4index_auto_in_arvalid),
    .auto_in_arid(axi4index_auto_in_arid),
    .auto_in_araddr(axi4index_auto_in_araddr),
    .auto_in_arlen(axi4index_auto_in_arlen),
    .auto_in_arsize(axi4index_auto_in_arsize),
    .auto_in_arburst(axi4index_auto_in_arburst),
    .auto_in_rready(axi4index_auto_in_rready),
    .auto_in_rvalid(axi4index_auto_in_rvalid),
    .auto_in_rid(axi4index_auto_in_rid),
    .auto_in_rdata(axi4index_auto_in_rdata),
    .auto_in_rresp(axi4index_auto_in_rresp),
    .auto_in_rlast(axi4index_auto_in_rlast),
    .auto_out_awready(axi4index_auto_out_awready),
    .auto_out_awvalid(axi4index_auto_out_awvalid),
    .auto_out_awid(axi4index_auto_out_awid),
    .auto_out_awaddr(axi4index_auto_out_awaddr),
    .auto_out_awlen(axi4index_auto_out_awlen),
    .auto_out_awsize(axi4index_auto_out_awsize),
    .auto_out_awburst(axi4index_auto_out_awburst),
    .auto_out_awecho_extra_id(axi4index_auto_out_awecho_extra_id),
    .auto_out_wready(axi4index_auto_out_wready),
    .auto_out_wvalid(axi4index_auto_out_wvalid),
    .auto_out_wdata(axi4index_auto_out_wdata),
    .auto_out_wstrb(axi4index_auto_out_wstrb),
    .auto_out_wlast(axi4index_auto_out_wlast),
    .auto_out_bready(axi4index_auto_out_bready),
    .auto_out_bvalid(axi4index_auto_out_bvalid),
    .auto_out_bid(axi4index_auto_out_bid),
    .auto_out_bresp(axi4index_auto_out_bresp),
    .auto_out_becho_extra_id(axi4index_auto_out_becho_extra_id),
    .auto_out_arready(axi4index_auto_out_arready),
    .auto_out_arvalid(axi4index_auto_out_arvalid),
    .auto_out_arid(axi4index_auto_out_arid),
    .auto_out_araddr(axi4index_auto_out_araddr),
    .auto_out_arlen(axi4index_auto_out_arlen),
    .auto_out_arsize(axi4index_auto_out_arsize),
    .auto_out_arburst(axi4index_auto_out_arburst),
    .auto_out_arecho_extra_id(axi4index_auto_out_arecho_extra_id),
    .auto_out_rready(axi4index_auto_out_rready),
    .auto_out_rvalid(axi4index_auto_out_rvalid),
    .auto_out_rid(axi4index_auto_out_rid),
    .auto_out_rdata(axi4index_auto_out_rdata),
    .auto_out_rresp(axi4index_auto_out_rresp),
    .auto_out_recho_extra_id(axi4index_auto_out_recho_extra_id),
    .auto_out_rlast(axi4index_auto_out_rlast)
  );
  AXI4UserYanker_1 axi4yank_1 ( // @[UserYanker.scala 105:30]
    .clock(axi4yank_1_clock),
    .reset(axi4yank_1_reset),
    .auto_in_awready(axi4yank_1_auto_in_awready),
    .auto_in_awvalid(axi4yank_1_auto_in_awvalid),
    .auto_in_awid(axi4yank_1_auto_in_awid),
    .auto_in_awaddr(axi4yank_1_auto_in_awaddr),
    .auto_in_awlen(axi4yank_1_auto_in_awlen),
    .auto_in_awsize(axi4yank_1_auto_in_awsize),
    .auto_in_awburst(axi4yank_1_auto_in_awburst),
    .auto_in_awecho_tl_state_size(axi4yank_1_auto_in_awecho_tl_state_size),
    .auto_in_awecho_tl_state_source(axi4yank_1_auto_in_awecho_tl_state_source),
    .auto_in_awecho_extra_id(axi4yank_1_auto_in_awecho_extra_id),
    .auto_in_wready(axi4yank_1_auto_in_wready),
    .auto_in_wvalid(axi4yank_1_auto_in_wvalid),
    .auto_in_wdata(axi4yank_1_auto_in_wdata),
    .auto_in_wstrb(axi4yank_1_auto_in_wstrb),
    .auto_in_wlast(axi4yank_1_auto_in_wlast),
    .auto_in_bready(axi4yank_1_auto_in_bready),
    .auto_in_bvalid(axi4yank_1_auto_in_bvalid),
    .auto_in_bid(axi4yank_1_auto_in_bid),
    .auto_in_bresp(axi4yank_1_auto_in_bresp),
    .auto_in_becho_tl_state_size(axi4yank_1_auto_in_becho_tl_state_size),
    .auto_in_becho_tl_state_source(axi4yank_1_auto_in_becho_tl_state_source),
    .auto_in_becho_extra_id(axi4yank_1_auto_in_becho_extra_id),
    .auto_in_arready(axi4yank_1_auto_in_arready),
    .auto_in_arvalid(axi4yank_1_auto_in_arvalid),
    .auto_in_arid(axi4yank_1_auto_in_arid),
    .auto_in_araddr(axi4yank_1_auto_in_araddr),
    .auto_in_arlen(axi4yank_1_auto_in_arlen),
    .auto_in_arsize(axi4yank_1_auto_in_arsize),
    .auto_in_arburst(axi4yank_1_auto_in_arburst),
    .auto_in_arecho_tl_state_size(axi4yank_1_auto_in_arecho_tl_state_size),
    .auto_in_arecho_tl_state_source(axi4yank_1_auto_in_arecho_tl_state_source),
    .auto_in_arecho_extra_id(axi4yank_1_auto_in_arecho_extra_id),
    .auto_in_rready(axi4yank_1_auto_in_rready),
    .auto_in_rvalid(axi4yank_1_auto_in_rvalid),
    .auto_in_rid(axi4yank_1_auto_in_rid),
    .auto_in_rdata(axi4yank_1_auto_in_rdata),
    .auto_in_rresp(axi4yank_1_auto_in_rresp),
    .auto_in_recho_tl_state_size(axi4yank_1_auto_in_recho_tl_state_size),
    .auto_in_recho_tl_state_source(axi4yank_1_auto_in_recho_tl_state_source),
    .auto_in_recho_extra_id(axi4yank_1_auto_in_recho_extra_id),
    .auto_in_rlast(axi4yank_1_auto_in_rlast),
    .auto_out_awready(axi4yank_1_auto_out_awready),
    .auto_out_awvalid(axi4yank_1_auto_out_awvalid),
    .auto_out_awid(axi4yank_1_auto_out_awid),
    .auto_out_awaddr(axi4yank_1_auto_out_awaddr),
    .auto_out_awlen(axi4yank_1_auto_out_awlen),
    .auto_out_awsize(axi4yank_1_auto_out_awsize),
    .auto_out_awburst(axi4yank_1_auto_out_awburst),
    .auto_out_wready(axi4yank_1_auto_out_wready),
    .auto_out_wvalid(axi4yank_1_auto_out_wvalid),
    .auto_out_wdata(axi4yank_1_auto_out_wdata),
    .auto_out_wstrb(axi4yank_1_auto_out_wstrb),
    .auto_out_wlast(axi4yank_1_auto_out_wlast),
    .auto_out_bready(axi4yank_1_auto_out_bready),
    .auto_out_bvalid(axi4yank_1_auto_out_bvalid),
    .auto_out_bid(axi4yank_1_auto_out_bid),
    .auto_out_bresp(axi4yank_1_auto_out_bresp),
    .auto_out_arready(axi4yank_1_auto_out_arready),
    .auto_out_arvalid(axi4yank_1_auto_out_arvalid),
    .auto_out_arid(axi4yank_1_auto_out_arid),
    .auto_out_araddr(axi4yank_1_auto_out_araddr),
    .auto_out_arlen(axi4yank_1_auto_out_arlen),
    .auto_out_arsize(axi4yank_1_auto_out_arsize),
    .auto_out_arburst(axi4yank_1_auto_out_arburst),
    .auto_out_rready(axi4yank_1_auto_out_rready),
    .auto_out_rvalid(axi4yank_1_auto_out_rvalid),
    .auto_out_rid(axi4yank_1_auto_out_rid),
    .auto_out_rdata(axi4yank_1_auto_out_rdata),
    .auto_out_rresp(axi4yank_1_auto_out_rresp),
    .auto_out_rlast(axi4yank_1_auto_out_rlast)
  );
  AXI4IdIndexer_1 axi4index_1 ( // @[IdIndexer.scala 91:31]
    .auto_in_awready(axi4index_1_auto_in_awready),
    .auto_in_awvalid(axi4index_1_auto_in_awvalid),
    .auto_in_awid(axi4index_1_auto_in_awid),
    .auto_in_awaddr(axi4index_1_auto_in_awaddr),
    .auto_in_awlen(axi4index_1_auto_in_awlen),
    .auto_in_awsize(axi4index_1_auto_in_awsize),
    .auto_in_awburst(axi4index_1_auto_in_awburst),
    .auto_in_awecho_tl_state_size(axi4index_1_auto_in_awecho_tl_state_size),
    .auto_in_awecho_tl_state_source(axi4index_1_auto_in_awecho_tl_state_source),
    .auto_in_wready(axi4index_1_auto_in_wready),
    .auto_in_wvalid(axi4index_1_auto_in_wvalid),
    .auto_in_wdata(axi4index_1_auto_in_wdata),
    .auto_in_wstrb(axi4index_1_auto_in_wstrb),
    .auto_in_wlast(axi4index_1_auto_in_wlast),
    .auto_in_bready(axi4index_1_auto_in_bready),
    .auto_in_bvalid(axi4index_1_auto_in_bvalid),
    .auto_in_bid(axi4index_1_auto_in_bid),
    .auto_in_bresp(axi4index_1_auto_in_bresp),
    .auto_in_becho_tl_state_size(axi4index_1_auto_in_becho_tl_state_size),
    .auto_in_becho_tl_state_source(axi4index_1_auto_in_becho_tl_state_source),
    .auto_in_arready(axi4index_1_auto_in_arready),
    .auto_in_arvalid(axi4index_1_auto_in_arvalid),
    .auto_in_arid(axi4index_1_auto_in_arid),
    .auto_in_araddr(axi4index_1_auto_in_araddr),
    .auto_in_arlen(axi4index_1_auto_in_arlen),
    .auto_in_arsize(axi4index_1_auto_in_arsize),
    .auto_in_arburst(axi4index_1_auto_in_arburst),
    .auto_in_arecho_tl_state_size(axi4index_1_auto_in_arecho_tl_state_size),
    .auto_in_arecho_tl_state_source(axi4index_1_auto_in_arecho_tl_state_source),
    .auto_in_rready(axi4index_1_auto_in_rready),
    .auto_in_rvalid(axi4index_1_auto_in_rvalid),
    .auto_in_rid(axi4index_1_auto_in_rid),
    .auto_in_rdata(axi4index_1_auto_in_rdata),
    .auto_in_rresp(axi4index_1_auto_in_rresp),
    .auto_in_recho_tl_state_size(axi4index_1_auto_in_recho_tl_state_size),
    .auto_in_recho_tl_state_source(axi4index_1_auto_in_recho_tl_state_source),
    .auto_in_rlast(axi4index_1_auto_in_rlast),
    .auto_out_awready(axi4index_1_auto_out_awready),
    .auto_out_awvalid(axi4index_1_auto_out_awvalid),
    .auto_out_awid(axi4index_1_auto_out_awid),
    .auto_out_awaddr(axi4index_1_auto_out_awaddr),
    .auto_out_awlen(axi4index_1_auto_out_awlen),
    .auto_out_awsize(axi4index_1_auto_out_awsize),
    .auto_out_awburst(axi4index_1_auto_out_awburst),
    .auto_out_awecho_tl_state_size(axi4index_1_auto_out_awecho_tl_state_size),
    .auto_out_awecho_tl_state_source(axi4index_1_auto_out_awecho_tl_state_source),
    .auto_out_awecho_extra_id(axi4index_1_auto_out_awecho_extra_id),
    .auto_out_wready(axi4index_1_auto_out_wready),
    .auto_out_wvalid(axi4index_1_auto_out_wvalid),
    .auto_out_wdata(axi4index_1_auto_out_wdata),
    .auto_out_wstrb(axi4index_1_auto_out_wstrb),
    .auto_out_wlast(axi4index_1_auto_out_wlast),
    .auto_out_bready(axi4index_1_auto_out_bready),
    .auto_out_bvalid(axi4index_1_auto_out_bvalid),
    .auto_out_bid(axi4index_1_auto_out_bid),
    .auto_out_bresp(axi4index_1_auto_out_bresp),
    .auto_out_becho_tl_state_size(axi4index_1_auto_out_becho_tl_state_size),
    .auto_out_becho_tl_state_source(axi4index_1_auto_out_becho_tl_state_source),
    .auto_out_becho_extra_id(axi4index_1_auto_out_becho_extra_id),
    .auto_out_arready(axi4index_1_auto_out_arready),
    .auto_out_arvalid(axi4index_1_auto_out_arvalid),
    .auto_out_arid(axi4index_1_auto_out_arid),
    .auto_out_araddr(axi4index_1_auto_out_araddr),
    .auto_out_arlen(axi4index_1_auto_out_arlen),
    .auto_out_arsize(axi4index_1_auto_out_arsize),
    .auto_out_arburst(axi4index_1_auto_out_arburst),
    .auto_out_arecho_tl_state_size(axi4index_1_auto_out_arecho_tl_state_size),
    .auto_out_arecho_tl_state_source(axi4index_1_auto_out_arecho_tl_state_source),
    .auto_out_arecho_extra_id(axi4index_1_auto_out_arecho_extra_id),
    .auto_out_rready(axi4index_1_auto_out_rready),
    .auto_out_rvalid(axi4index_1_auto_out_rvalid),
    .auto_out_rid(axi4index_1_auto_out_rid),
    .auto_out_rdata(axi4index_1_auto_out_rdata),
    .auto_out_rresp(axi4index_1_auto_out_rresp),
    .auto_out_recho_tl_state_size(axi4index_1_auto_out_recho_tl_state_size),
    .auto_out_recho_tl_state_source(axi4index_1_auto_out_recho_tl_state_source),
    .auto_out_recho_extra_id(axi4index_1_auto_out_recho_extra_id),
    .auto_out_rlast(axi4index_1_auto_out_rlast)
  );
  TLToAXI4 tl2axi4 ( // @[ToAXI4.scala 283:29]
    .clock(tl2axi4_clock),
    .reset(tl2axi4_reset),
    .auto_in_a_ready(tl2axi4_auto_in_a_ready),
    .auto_in_a_valid(tl2axi4_auto_in_a_valid),
    .auto_in_a_bits_opcode(tl2axi4_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(tl2axi4_auto_in_a_bits_param),
    .auto_in_a_bits_size(tl2axi4_auto_in_a_bits_size),
    .auto_in_a_bits_source(tl2axi4_auto_in_a_bits_source),
    .auto_in_a_bits_address(tl2axi4_auto_in_a_bits_address),
    .auto_in_a_bits_mask(tl2axi4_auto_in_a_bits_mask),
    .auto_in_a_bits_data(tl2axi4_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(tl2axi4_auto_in_a_bits_corrupt),
    .auto_in_d_ready(tl2axi4_auto_in_d_ready),
    .auto_in_d_valid(tl2axi4_auto_in_d_valid),
    .auto_in_d_bits_opcode(tl2axi4_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(tl2axi4_auto_in_d_bits_size),
    .auto_in_d_bits_source(tl2axi4_auto_in_d_bits_source),
    .auto_in_d_bits_denied(tl2axi4_auto_in_d_bits_denied),
    .auto_in_d_bits_data(tl2axi4_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(tl2axi4_auto_in_d_bits_corrupt),
    .auto_out_awready(tl2axi4_auto_out_awready),
    .auto_out_awvalid(tl2axi4_auto_out_awvalid),
    .auto_out_awid(tl2axi4_auto_out_awid),
    .auto_out_awaddr(tl2axi4_auto_out_awaddr),
    .auto_out_awlen(tl2axi4_auto_out_awlen),
    .auto_out_awsize(tl2axi4_auto_out_awsize),
    .auto_out_awburst(tl2axi4_auto_out_awburst),
    .auto_out_awecho_tl_state_size(tl2axi4_auto_out_awecho_tl_state_size),
    .auto_out_awecho_tl_state_source(tl2axi4_auto_out_awecho_tl_state_source),
    .auto_out_wready(tl2axi4_auto_out_wready),
    .auto_out_wvalid(tl2axi4_auto_out_wvalid),
    .auto_out_wdata(tl2axi4_auto_out_wdata),
    .auto_out_wstrb(tl2axi4_auto_out_wstrb),
    .auto_out_wlast(tl2axi4_auto_out_wlast),
    .auto_out_bready(tl2axi4_auto_out_bready),
    .auto_out_bvalid(tl2axi4_auto_out_bvalid),
    .auto_out_bid(tl2axi4_auto_out_bid),
    .auto_out_bresp(tl2axi4_auto_out_bresp),
    .auto_out_becho_tl_state_size(tl2axi4_auto_out_becho_tl_state_size),
    .auto_out_becho_tl_state_source(tl2axi4_auto_out_becho_tl_state_source),
    .auto_out_arready(tl2axi4_auto_out_arready),
    .auto_out_arvalid(tl2axi4_auto_out_arvalid),
    .auto_out_arid(tl2axi4_auto_out_arid),
    .auto_out_araddr(tl2axi4_auto_out_araddr),
    .auto_out_arlen(tl2axi4_auto_out_arlen),
    .auto_out_arsize(tl2axi4_auto_out_arsize),
    .auto_out_arburst(tl2axi4_auto_out_arburst),
    .auto_out_arecho_tl_state_size(tl2axi4_auto_out_arecho_tl_state_size),
    .auto_out_arecho_tl_state_source(tl2axi4_auto_out_arecho_tl_state_source),
    .auto_out_rready(tl2axi4_auto_out_rready),
    .auto_out_rvalid(tl2axi4_auto_out_rvalid),
    .auto_out_rid(tl2axi4_auto_out_rid),
    .auto_out_rdata(tl2axi4_auto_out_rdata),
    .auto_out_rresp(tl2axi4_auto_out_rresp),
    .auto_out_recho_tl_state_size(tl2axi4_auto_out_recho_tl_state_size),
    .auto_out_recho_tl_state_source(tl2axi4_auto_out_recho_tl_state_source),
    .auto_out_rlast(tl2axi4_auto_out_rlast)
  );
  TLError_2 err ( // @[ChipLinkBridge.scala 150:23]
    .clock(err_clock),
    .reset(err_reset),
    .auto_in_a_ready(err_auto_in_a_ready),
    .auto_in_a_valid(err_auto_in_a_valid),
    .auto_in_a_bits_opcode(err_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(err_auto_in_a_bits_param),
    .auto_in_a_bits_size(err_auto_in_a_bits_size),
    .auto_in_a_bits_source(err_auto_in_a_bits_source),
    .auto_in_a_bits_address(err_auto_in_a_bits_address),
    .auto_in_a_bits_mask(err_auto_in_a_bits_mask),
    .auto_in_a_bits_corrupt(err_auto_in_a_bits_corrupt),
    .auto_in_c_ready(err_auto_in_c_ready),
    .auto_in_c_valid(err_auto_in_c_valid),
    .auto_in_c_bits_opcode(err_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(err_auto_in_c_bits_param),
    .auto_in_c_bits_size(err_auto_in_c_bits_size),
    .auto_in_c_bits_source(err_auto_in_c_bits_source),
    .auto_in_c_bits_address(err_auto_in_c_bits_address),
    .auto_in_d_ready(err_auto_in_d_ready),
    .auto_in_d_valid(err_auto_in_d_valid),
    .auto_in_d_bits_opcode(err_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(err_auto_in_d_bits_param),
    .auto_in_d_bits_size(err_auto_in_d_bits_size),
    .auto_in_d_bits_source(err_auto_in_d_bits_source),
    .auto_in_d_bits_denied(err_auto_in_d_bits_denied),
    .auto_in_d_bits_corrupt(err_auto_in_d_bits_corrupt),
    .auto_in_e_valid(err_auto_in_e_valid)
  );
  TLAtomicAutomata atomics ( // @[AtomicAutomata.scala 283:29]
    .clock(atomics_clock),
    .reset(atomics_reset),
    .auto_in_a_ready(atomics_auto_in_a_ready),
    .auto_in_a_valid(atomics_auto_in_a_valid),
    .auto_in_a_bits_opcode(atomics_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(atomics_auto_in_a_bits_param),
    .auto_in_a_bits_size(atomics_auto_in_a_bits_size),
    .auto_in_a_bits_source(atomics_auto_in_a_bits_source),
    .auto_in_a_bits_address(atomics_auto_in_a_bits_address),
    .auto_in_a_bits_mask(atomics_auto_in_a_bits_mask),
    .auto_in_a_bits_data(atomics_auto_in_a_bits_data),
    .auto_in_c_ready(atomics_auto_in_c_ready),
    .auto_in_c_valid(atomics_auto_in_c_valid),
    .auto_in_c_bits_opcode(atomics_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(atomics_auto_in_c_bits_param),
    .auto_in_c_bits_size(atomics_auto_in_c_bits_size),
    .auto_in_c_bits_source(atomics_auto_in_c_bits_source),
    .auto_in_c_bits_address(atomics_auto_in_c_bits_address),
    .auto_in_d_ready(atomics_auto_in_d_ready),
    .auto_in_d_valid(atomics_auto_in_d_valid),
    .auto_in_d_bits_opcode(atomics_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(atomics_auto_in_d_bits_param),
    .auto_in_d_bits_size(atomics_auto_in_d_bits_size),
    .auto_in_d_bits_source(atomics_auto_in_d_bits_source),
    .auto_in_d_bits_denied(atomics_auto_in_d_bits_denied),
    .auto_in_d_bits_data(atomics_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(atomics_auto_in_d_bits_corrupt),
    .auto_in_e_ready(atomics_auto_in_e_ready),
    .auto_in_e_valid(atomics_auto_in_e_valid),
    .auto_in_e_bits_sink(atomics_auto_in_e_bits_sink),
    .auto_out_a_ready(atomics_auto_out_a_ready),
    .auto_out_a_valid(atomics_auto_out_a_valid),
    .auto_out_a_bits_opcode(atomics_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(atomics_auto_out_a_bits_param),
    .auto_out_a_bits_size(atomics_auto_out_a_bits_size),
    .auto_out_a_bits_source(atomics_auto_out_a_bits_source),
    .auto_out_a_bits_address(atomics_auto_out_a_bits_address),
    .auto_out_a_bits_mask(atomics_auto_out_a_bits_mask),
    .auto_out_a_bits_data(atomics_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(atomics_auto_out_a_bits_corrupt),
    .auto_out_c_ready(atomics_auto_out_c_ready),
    .auto_out_c_valid(atomics_auto_out_c_valid),
    .auto_out_c_bits_opcode(atomics_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(atomics_auto_out_c_bits_param),
    .auto_out_c_bits_size(atomics_auto_out_c_bits_size),
    .auto_out_c_bits_source(atomics_auto_out_c_bits_source),
    .auto_out_c_bits_address(atomics_auto_out_c_bits_address),
    .auto_out_d_ready(atomics_auto_out_d_ready),
    .auto_out_d_valid(atomics_auto_out_d_valid),
    .auto_out_d_bits_opcode(atomics_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(atomics_auto_out_d_bits_param),
    .auto_out_d_bits_size(atomics_auto_out_d_bits_size),
    .auto_out_d_bits_source(atomics_auto_out_d_bits_source),
    .auto_out_d_bits_denied(atomics_auto_out_d_bits_denied),
    .auto_out_d_bits_data(atomics_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(atomics_auto_out_d_bits_corrupt),
    .auto_out_e_ready(atomics_auto_out_e_ready),
    .auto_out_e_valid(atomics_auto_out_e_valid),
    .auto_out_e_bits_sink(atomics_auto_out_e_bits_sink)
  );
  TLFIFOFixer_1 fixer_1 ( // @[FIFOFixer.scala 144:27]
    .clock(fixer_1_clock),
    .reset(fixer_1_reset),
    .auto_in_a_ready(fixer_1_auto_in_a_ready),
    .auto_in_a_valid(fixer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fixer_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(fixer_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_1_auto_in_a_bits_data),
    .auto_in_c_ready(fixer_1_auto_in_c_ready),
    .auto_in_c_valid(fixer_1_auto_in_c_valid),
    .auto_in_c_bits_opcode(fixer_1_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(fixer_1_auto_in_c_bits_param),
    .auto_in_c_bits_size(fixer_1_auto_in_c_bits_size),
    .auto_in_c_bits_source(fixer_1_auto_in_c_bits_source),
    .auto_in_c_bits_address(fixer_1_auto_in_c_bits_address),
    .auto_in_d_ready(fixer_1_auto_in_d_ready),
    .auto_in_d_valid(fixer_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fixer_1_auto_in_d_bits_param),
    .auto_in_d_bits_size(fixer_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_1_auto_in_d_bits_source),
    .auto_in_d_bits_denied(fixer_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_1_auto_in_d_bits_corrupt),
    .auto_in_e_ready(fixer_1_auto_in_e_ready),
    .auto_in_e_valid(fixer_1_auto_in_e_valid),
    .auto_in_e_bits_sink(fixer_1_auto_in_e_bits_sink),
    .auto_out_a_ready(fixer_1_auto_out_a_ready),
    .auto_out_a_valid(fixer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fixer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(fixer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_1_auto_out_a_bits_data),
    .auto_out_c_ready(fixer_1_auto_out_c_ready),
    .auto_out_c_valid(fixer_1_auto_out_c_valid),
    .auto_out_c_bits_opcode(fixer_1_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(fixer_1_auto_out_c_bits_param),
    .auto_out_c_bits_size(fixer_1_auto_out_c_bits_size),
    .auto_out_c_bits_source(fixer_1_auto_out_c_bits_source),
    .auto_out_c_bits_address(fixer_1_auto_out_c_bits_address),
    .auto_out_d_ready(fixer_1_auto_out_d_ready),
    .auto_out_d_valid(fixer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fixer_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(fixer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_1_auto_out_d_bits_source),
    .auto_out_d_bits_denied(fixer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_1_auto_out_d_bits_corrupt),
    .auto_out_e_ready(fixer_1_auto_out_e_ready),
    .auto_out_e_valid(fixer_1_auto_out_e_valid),
    .auto_out_e_bits_sink(fixer_1_auto_out_e_bits_sink)
  );
  TLHintHandler hints ( // @[HintHandler.scala 119:27]
    .clock(hints_clock),
    .reset(hints_reset),
    .auto_in_a_ready(hints_auto_in_a_ready),
    .auto_in_a_valid(hints_auto_in_a_valid),
    .auto_in_a_bits_opcode(hints_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(hints_auto_in_a_bits_param),
    .auto_in_a_bits_size(hints_auto_in_a_bits_size),
    .auto_in_a_bits_source(hints_auto_in_a_bits_source),
    .auto_in_a_bits_address(hints_auto_in_a_bits_address),
    .auto_in_a_bits_mask(hints_auto_in_a_bits_mask),
    .auto_in_a_bits_data(hints_auto_in_a_bits_data),
    .auto_in_c_ready(hints_auto_in_c_ready),
    .auto_in_c_valid(hints_auto_in_c_valid),
    .auto_in_c_bits_opcode(hints_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(hints_auto_in_c_bits_param),
    .auto_in_c_bits_size(hints_auto_in_c_bits_size),
    .auto_in_c_bits_source(hints_auto_in_c_bits_source),
    .auto_in_c_bits_address(hints_auto_in_c_bits_address),
    .auto_in_d_ready(hints_auto_in_d_ready),
    .auto_in_d_valid(hints_auto_in_d_valid),
    .auto_in_d_bits_opcode(hints_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(hints_auto_in_d_bits_param),
    .auto_in_d_bits_size(hints_auto_in_d_bits_size),
    .auto_in_d_bits_source(hints_auto_in_d_bits_source),
    .auto_in_d_bits_denied(hints_auto_in_d_bits_denied),
    .auto_in_d_bits_data(hints_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(hints_auto_in_d_bits_corrupt),
    .auto_in_e_ready(hints_auto_in_e_ready),
    .auto_in_e_valid(hints_auto_in_e_valid),
    .auto_in_e_bits_sink(hints_auto_in_e_bits_sink),
    .auto_out_a_ready(hints_auto_out_a_ready),
    .auto_out_a_valid(hints_auto_out_a_valid),
    .auto_out_a_bits_opcode(hints_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(hints_auto_out_a_bits_param),
    .auto_out_a_bits_size(hints_auto_out_a_bits_size),
    .auto_out_a_bits_source(hints_auto_out_a_bits_source),
    .auto_out_a_bits_address(hints_auto_out_a_bits_address),
    .auto_out_a_bits_mask(hints_auto_out_a_bits_mask),
    .auto_out_a_bits_data(hints_auto_out_a_bits_data),
    .auto_out_c_ready(hints_auto_out_c_ready),
    .auto_out_c_valid(hints_auto_out_c_valid),
    .auto_out_c_bits_opcode(hints_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(hints_auto_out_c_bits_param),
    .auto_out_c_bits_size(hints_auto_out_c_bits_size),
    .auto_out_c_bits_source(hints_auto_out_c_bits_source),
    .auto_out_c_bits_address(hints_auto_out_c_bits_address),
    .auto_out_d_ready(hints_auto_out_d_ready),
    .auto_out_d_valid(hints_auto_out_d_valid),
    .auto_out_d_bits_opcode(hints_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(hints_auto_out_d_bits_param),
    .auto_out_d_bits_size(hints_auto_out_d_bits_size),
    .auto_out_d_bits_source(hints_auto_out_d_bits_source),
    .auto_out_d_bits_denied(hints_auto_out_d_bits_denied),
    .auto_out_d_bits_data(hints_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(hints_auto_out_d_bits_corrupt),
    .auto_out_e_ready(hints_auto_out_e_ready),
    .auto_out_e_valid(hints_auto_out_e_valid),
    .auto_out_e_bits_sink(hints_auto_out_e_bits_sink)
  );
  TLWidthWidget_1 widget_1 ( // @[WidthWidget.scala 219:28]
    .clock(widget_1_clock),
    .reset(widget_1_reset),
    .auto_in_a_ready(widget_1_auto_in_a_ready),
    .auto_in_a_valid(widget_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(widget_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(widget_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_1_auto_in_a_bits_data),
    .auto_in_c_ready(widget_1_auto_in_c_ready),
    .auto_in_c_valid(widget_1_auto_in_c_valid),
    .auto_in_c_bits_opcode(widget_1_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(widget_1_auto_in_c_bits_param),
    .auto_in_c_bits_size(widget_1_auto_in_c_bits_size),
    .auto_in_c_bits_source(widget_1_auto_in_c_bits_source),
    .auto_in_c_bits_address(widget_1_auto_in_c_bits_address),
    .auto_in_d_ready(widget_1_auto_in_d_ready),
    .auto_in_d_valid(widget_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(widget_1_auto_in_d_bits_param),
    .auto_in_d_bits_size(widget_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_1_auto_in_d_bits_source),
    .auto_in_d_bits_denied(widget_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_1_auto_in_d_bits_corrupt),
    .auto_in_e_ready(widget_1_auto_in_e_ready),
    .auto_in_e_valid(widget_1_auto_in_e_valid),
    .auto_in_e_bits_sink(widget_1_auto_in_e_bits_sink),
    .auto_out_a_ready(widget_1_auto_out_a_ready),
    .auto_out_a_valid(widget_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(widget_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(widget_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_1_auto_out_a_bits_data),
    .auto_out_c_ready(widget_1_auto_out_c_ready),
    .auto_out_c_valid(widget_1_auto_out_c_valid),
    .auto_out_c_bits_opcode(widget_1_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(widget_1_auto_out_c_bits_param),
    .auto_out_c_bits_size(widget_1_auto_out_c_bits_size),
    .auto_out_c_bits_source(widget_1_auto_out_c_bits_source),
    .auto_out_c_bits_address(widget_1_auto_out_c_bits_address),
    .auto_out_d_ready(widget_1_auto_out_d_ready),
    .auto_out_d_valid(widget_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_1_auto_out_d_bits_source),
    .auto_out_d_bits_denied(widget_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_1_auto_out_d_bits_corrupt),
    .auto_out_e_ready(widget_1_auto_out_e_ready),
    .auto_out_e_valid(widget_1_auto_out_e_valid),
    .auto_out_e_bits_sink(widget_1_auto_out_e_bits_sink)
  );
  TLWidthWidget_2 widget_2 ( // @[WidthWidget.scala 219:28]
    .clock(widget_2_clock),
    .reset(widget_2_reset),
    .auto_in_a_ready(widget_2_auto_in_a_ready),
    .auto_in_a_valid(widget_2_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_2_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(widget_2_auto_in_a_bits_param),
    .auto_in_a_bits_size(widget_2_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_2_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_2_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_2_auto_in_a_bits_mask),
    .auto_in_a_bits_corrupt(widget_2_auto_in_a_bits_corrupt),
    .auto_in_c_ready(widget_2_auto_in_c_ready),
    .auto_in_c_valid(widget_2_auto_in_c_valid),
    .auto_in_c_bits_opcode(widget_2_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(widget_2_auto_in_c_bits_param),
    .auto_in_c_bits_size(widget_2_auto_in_c_bits_size),
    .auto_in_c_bits_source(widget_2_auto_in_c_bits_source),
    .auto_in_c_bits_address(widget_2_auto_in_c_bits_address),
    .auto_in_d_ready(widget_2_auto_in_d_ready),
    .auto_in_d_valid(widget_2_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_2_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(widget_2_auto_in_d_bits_param),
    .auto_in_d_bits_size(widget_2_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_2_auto_in_d_bits_source),
    .auto_in_d_bits_denied(widget_2_auto_in_d_bits_denied),
    .auto_in_d_bits_corrupt(widget_2_auto_in_d_bits_corrupt),
    .auto_in_e_valid(widget_2_auto_in_e_valid),
    .auto_out_a_ready(widget_2_auto_out_a_ready),
    .auto_out_a_valid(widget_2_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_2_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(widget_2_auto_out_a_bits_param),
    .auto_out_a_bits_size(widget_2_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_2_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_2_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_2_auto_out_a_bits_mask),
    .auto_out_a_bits_corrupt(widget_2_auto_out_a_bits_corrupt),
    .auto_out_c_ready(widget_2_auto_out_c_ready),
    .auto_out_c_valid(widget_2_auto_out_c_valid),
    .auto_out_c_bits_opcode(widget_2_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(widget_2_auto_out_c_bits_param),
    .auto_out_c_bits_size(widget_2_auto_out_c_bits_size),
    .auto_out_c_bits_source(widget_2_auto_out_c_bits_source),
    .auto_out_c_bits_address(widget_2_auto_out_c_bits_address),
    .auto_out_d_ready(widget_2_auto_out_d_ready),
    .auto_out_d_valid(widget_2_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_2_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_2_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_2_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_2_auto_out_d_bits_source),
    .auto_out_d_bits_denied(widget_2_auto_out_d_bits_denied),
    .auto_out_d_bits_corrupt(widget_2_auto_out_d_bits_corrupt),
    .auto_out_e_valid(widget_2_auto_out_e_valid)
  );
  assign slave_0_awready = axi4index_auto_in_awready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_wready = axi4index_auto_in_wready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_bvalid = axi4index_auto_in_bvalid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_bid = axi4index_auto_in_bid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_bresp = axi4index_auto_in_bresp; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_arready = axi4index_auto_in_arready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_rvalid = axi4index_auto_in_rvalid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_rid = axi4index_auto_in_rid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_rdata = axi4index_auto_in_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_rresp = axi4index_auto_in_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign slave_0_rlast = axi4index_auto_in_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign master_mem_0_awvalid = axi4yank_1_auto_out_awvalid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_awid = axi4yank_1_auto_out_awid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_awaddr = axi4yank_1_auto_out_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_awlen = axi4yank_1_auto_out_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_awsize = axi4yank_1_auto_out_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_awburst = axi4yank_1_auto_out_awburst; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_wvalid = axi4yank_1_auto_out_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_wdata = axi4yank_1_auto_out_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_wstrb = axi4yank_1_auto_out_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_wlast = axi4yank_1_auto_out_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_bready = axi4yank_1_auto_out_bready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_arvalid = axi4yank_1_auto_out_arvalid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_arid = axi4yank_1_auto_out_arid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_araddr = axi4yank_1_auto_out_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_arlen = axi4yank_1_auto_out_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_arsize = axi4yank_1_auto_out_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_arburst = axi4yank_1_auto_out_arburst; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign master_mem_0_rready = axi4yank_1_auto_out_rready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign fpga_io_c2b_clk = chiplink_auto_io_out_c2b_clk; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign fpga_io_c2b_rst = chiplink_auto_io_out_c2b_rst; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign fpga_io_c2b_send = chiplink_auto_io_out_c2b_send; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign fpga_io_c2b_data = chiplink_auto_io_out_c2b_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_auto_in_a_valid = atomics_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_a_bits_opcode = atomics_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_a_bits_param = atomics_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_a_bits_size = atomics_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_a_bits_source = atomics_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_a_bits_address = atomics_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_a_bits_mask = atomics_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_a_bits_data = atomics_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_a_bits_corrupt = atomics_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_c_valid = atomics_auto_out_c_valid; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_c_bits_opcode = atomics_auto_out_c_bits_opcode; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_c_bits_param = atomics_auto_out_c_bits_param; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_c_bits_size = atomics_auto_out_c_bits_size; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_c_bits_source = atomics_auto_out_c_bits_source; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_c_bits_address = atomics_auto_out_c_bits_address; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_d_ready = atomics_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_e_valid = atomics_auto_out_e_valid; // @[LazyModule.scala 296:16]
  assign xbar_auto_in_e_bits_sink = atomics_auto_out_e_bits_sink; // @[LazyModule.scala 296:16]
  assign xbar_auto_out_1_a_ready = widget_2_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_1_c_ready = widget_2_auto_in_c_ready; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_1_d_valid = widget_2_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_1_d_bits_opcode = widget_2_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_1_d_bits_param = widget_2_auto_in_d_bits_param; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_1_d_bits_size = widget_2_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_1_d_bits_source = widget_2_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_1_d_bits_denied = widget_2_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_1_d_bits_corrupt = widget_2_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_0_a_ready = tl2axi4_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_0_d_valid = tl2axi4_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_0_d_bits_opcode = tl2axi4_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_0_d_bits_size = tl2axi4_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_0_d_bits_source = tl2axi4_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_0_d_bits_denied = tl2axi4_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_0_d_bits_data = tl2axi4_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign xbar_auto_out_0_d_bits_corrupt = tl2axi4_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign xbar_1_clock = clock;
  assign xbar_1_reset = reset;
  assign xbar_1_auto_in_a_valid = fixer_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_in_a_bits_data = fixer_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_in_d_ready = fixer_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_out_1_a_ready = ferr_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_1_d_valid = ferr_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_1_d_bits_opcode = ferr_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_1_d_bits_size = ferr_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_1_d_bits_source = ferr_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_1_d_bits_denied = ferr_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_1_d_bits_corrupt = ferr_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_a_ready = chiplink_auto_sbypass_node_in_in_a_ready; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_valid = chiplink_auto_sbypass_node_in_in_d_valid; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_bits_opcode = chiplink_auto_sbypass_node_in_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_bits_param = chiplink_auto_sbypass_node_in_in_d_bits_param; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_bits_size = chiplink_auto_sbypass_node_in_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_bits_source = chiplink_auto_sbypass_node_in_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_bits_sink = chiplink_auto_sbypass_node_in_in_d_bits_sink; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_bits_denied = chiplink_auto_sbypass_node_in_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_bits_data = chiplink_auto_sbypass_node_in_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign xbar_1_auto_out_0_d_bits_corrupt = chiplink_auto_sbypass_node_in_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign ferr_clock = clock;
  assign ferr_reset = reset;
  assign ferr_auto_in_a_valid = xbar_1_auto_out_1_a_valid; // @[LazyModule.scala 298:16]
  assign ferr_auto_in_a_bits_opcode = xbar_1_auto_out_1_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign ferr_auto_in_a_bits_size = xbar_1_auto_out_1_a_bits_size; // @[LazyModule.scala 298:16]
  assign ferr_auto_in_a_bits_source = xbar_1_auto_out_1_a_bits_source; // @[LazyModule.scala 298:16]
  assign ferr_auto_in_a_bits_address = xbar_1_auto_out_1_a_bits_address; // @[LazyModule.scala 298:16]
  assign ferr_auto_in_a_bits_mask = xbar_1_auto_out_1_a_bits_mask; // @[LazyModule.scala 298:16]
  assign ferr_auto_in_d_ready = xbar_1_auto_out_1_d_ready; // @[LazyModule.scala 298:16]
  assign chiplink_clock = clock;
  assign chiplink_reset = reset;
  assign chiplink_auto_mbypass_out_a_ready = widget_1_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_c_ready = widget_1_auto_in_c_ready; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_d_valid = widget_1_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_d_bits_opcode = widget_1_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_d_bits_param = widget_1_auto_in_d_bits_param; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_d_bits_size = widget_1_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_d_bits_source = widget_1_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_d_bits_denied = widget_1_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_d_bits_data = widget_1_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_d_bits_corrupt = widget_1_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign chiplink_auto_mbypass_out_e_ready = widget_1_auto_in_e_ready; // @[LazyModule.scala 298:16]
  assign chiplink_auto_sbypass_node_in_in_a_valid = xbar_1_auto_out_0_a_valid; // @[LazyModule.scala 298:16]
  assign chiplink_auto_sbypass_node_in_in_a_bits_opcode = xbar_1_auto_out_0_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign chiplink_auto_sbypass_node_in_in_a_bits_size = xbar_1_auto_out_0_a_bits_size; // @[LazyModule.scala 298:16]
  assign chiplink_auto_sbypass_node_in_in_a_bits_source = xbar_1_auto_out_0_a_bits_source; // @[LazyModule.scala 298:16]
  assign chiplink_auto_sbypass_node_in_in_a_bits_address = xbar_1_auto_out_0_a_bits_address; // @[LazyModule.scala 298:16]
  assign chiplink_auto_sbypass_node_in_in_a_bits_mask = xbar_1_auto_out_0_a_bits_mask; // @[LazyModule.scala 298:16]
  assign chiplink_auto_sbypass_node_in_in_a_bits_data = xbar_1_auto_out_0_a_bits_data; // @[LazyModule.scala 298:16]
  assign chiplink_auto_sbypass_node_in_in_d_ready = xbar_1_auto_out_0_d_ready; // @[LazyModule.scala 298:16]
  assign chiplink_auto_io_out_b2c_clk = fpga_io_b2c_clk; // @[Nodes.scala 1210:84 BundleBridge.scala 54:8]
  assign chiplink_auto_io_out_b2c_rst = fpga_io_b2c_rst; // @[Nodes.scala 1210:84 BundleBridge.scala 54:8]
  assign chiplink_auto_io_out_b2c_send = fpga_io_b2c_send; // @[Nodes.scala 1210:84 BundleBridge.scala 54:8]
  assign chiplink_auto_io_out_b2c_data = fpga_io_b2c_data; // @[Nodes.scala 1210:84 BundleBridge.scala 54:8]
  assign fixer_clock = clock;
  assign fixer_reset = reset;
  assign fixer_auto_in_a_valid = widget_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_size = widget_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_source = widget_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_address = widget_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_mask = widget_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_data = widget_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_d_ready = widget_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_a_ready = xbar_1_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_valid = xbar_1_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_opcode = xbar_1_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_param = xbar_1_auto_in_d_bits_param; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_size = xbar_1_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_source = xbar_1_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_sink = xbar_1_auto_in_d_bits_sink; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_denied = xbar_1_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_data = xbar_1_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_corrupt = xbar_1_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = axi42tl_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_opcode = axi42tl_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_size = axi42tl_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_source = axi42tl_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_address = axi42tl_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_mask = axi42tl_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_data = axi42tl_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign widget_auto_in_d_ready = axi42tl_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign widget_auto_out_a_ready = fixer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_valid = fixer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_param = fixer_auto_in_d_bits_param; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_size = fixer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_source = fixer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_sink = fixer_auto_in_d_bits_sink; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_data = fixer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign axi42tl_clock = clock;
  assign axi42tl_reset = reset;
  assign axi42tl_auto_in_awvalid = axi4yank_auto_out_awvalid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_awid = axi4yank_auto_out_awid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_awaddr = axi4yank_auto_out_awaddr; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_awlen = axi4yank_auto_out_awlen; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_awsize = axi4yank_auto_out_awsize; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_wvalid = axi4yank_auto_out_wvalid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_wdata = axi4yank_auto_out_wdata; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_wstrb = axi4yank_auto_out_wstrb; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_wlast = axi4yank_auto_out_wlast; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_bready = axi4yank_auto_out_bready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_arvalid = axi4yank_auto_out_arvalid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_arid = axi4yank_auto_out_arid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_araddr = axi4yank_auto_out_araddr; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_arlen = axi4yank_auto_out_arlen; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_arsize = axi4yank_auto_out_arsize; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_rready = axi4yank_auto_out_rready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_a_ready = widget_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_valid = widget_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_size = widget_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_source = widget_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_denied = widget_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_data = widget_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_corrupt = widget_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign axi4yank_clock = clock;
  assign axi4yank_reset = reset;
  assign axi4yank_auto_in_awvalid = axi4frag_auto_out_awvalid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_awid = axi4frag_auto_out_awid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_awaddr = axi4frag_auto_out_awaddr; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_awlen = axi4frag_auto_out_awlen; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_awsize = axi4frag_auto_out_awsize; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_awecho_extra_id = axi4frag_auto_out_awecho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_awecho_real_last = axi4frag_auto_out_awecho_real_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_wvalid = axi4frag_auto_out_wvalid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_wdata = axi4frag_auto_out_wdata; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_wstrb = axi4frag_auto_out_wstrb; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_wlast = axi4frag_auto_out_wlast; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_bready = axi4frag_auto_out_bready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_arvalid = axi4frag_auto_out_arvalid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_arid = axi4frag_auto_out_arid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_araddr = axi4frag_auto_out_araddr; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_arlen = axi4frag_auto_out_arlen; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_arsize = axi4frag_auto_out_arsize; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_arecho_extra_id = axi4frag_auto_out_arecho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_arecho_real_last = axi4frag_auto_out_arecho_real_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_rready = axi4frag_auto_out_rready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_awready = axi42tl_auto_in_awready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_wready = axi42tl_auto_in_wready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_bvalid = axi42tl_auto_in_bvalid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_bid = axi42tl_auto_in_bid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_bresp = axi42tl_auto_in_bresp; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_arready = axi42tl_auto_in_arready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_rvalid = axi42tl_auto_in_rvalid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_rid = axi42tl_auto_in_rid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_rdata = axi42tl_auto_in_rdata; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_rresp = axi42tl_auto_in_rresp; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_rlast = axi42tl_auto_in_rlast; // @[LazyModule.scala 296:16]
  assign axi4frag_clock = clock;
  assign axi4frag_reset = reset;
  assign axi4frag_auto_in_awvalid = axi4index_auto_out_awvalid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_awid = axi4index_auto_out_awid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_awaddr = axi4index_auto_out_awaddr; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_awlen = axi4index_auto_out_awlen; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_awsize = axi4index_auto_out_awsize; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_awburst = axi4index_auto_out_awburst; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_awecho_extra_id = axi4index_auto_out_awecho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_wvalid = axi4index_auto_out_wvalid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_wdata = axi4index_auto_out_wdata; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_wstrb = axi4index_auto_out_wstrb; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_wlast = axi4index_auto_out_wlast; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_bready = axi4index_auto_out_bready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_arvalid = axi4index_auto_out_arvalid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_arid = axi4index_auto_out_arid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_araddr = axi4index_auto_out_araddr; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_arlen = axi4index_auto_out_arlen; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_arsize = axi4index_auto_out_arsize; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_arburst = axi4index_auto_out_arburst; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_arecho_extra_id = axi4index_auto_out_arecho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_rready = axi4index_auto_out_rready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_awready = axi4yank_auto_in_awready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_wready = axi4yank_auto_in_wready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_bvalid = axi4yank_auto_in_bvalid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_bid = axi4yank_auto_in_bid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_bresp = axi4yank_auto_in_bresp; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_becho_extra_id = axi4yank_auto_in_becho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_becho_real_last = axi4yank_auto_in_becho_real_last; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_arready = axi4yank_auto_in_arready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_rvalid = axi4yank_auto_in_rvalid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_rid = axi4yank_auto_in_rid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_rdata = axi4yank_auto_in_rdata; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_rresp = axi4yank_auto_in_rresp; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_recho_extra_id = axi4yank_auto_in_recho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_recho_real_last = axi4yank_auto_in_recho_real_last; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_rlast = axi4yank_auto_in_rlast; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_awvalid = slave_0_awvalid; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_awid = slave_0_awid; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_awaddr = slave_0_awaddr; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_awlen = slave_0_awlen; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_awsize = slave_0_awsize; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_awburst = slave_0_awburst; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_wvalid = slave_0_wvalid; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_wdata = slave_0_wdata; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_wstrb = slave_0_wstrb; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_wlast = slave_0_wlast; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_bready = slave_0_bready; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_arvalid = slave_0_arvalid; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_arid = slave_0_arid; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_araddr = slave_0_araddr; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_arlen = slave_0_arlen; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_arsize = slave_0_arsize; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_arburst = slave_0_arburst; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_in_rready = slave_0_rready; // @[Nodes.scala 1207:84 Nodes.scala 1630:60]
  assign axi4index_auto_out_awready = axi4frag_auto_in_awready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_wready = axi4frag_auto_in_wready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_bvalid = axi4frag_auto_in_bvalid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_bid = axi4frag_auto_in_bid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_bresp = axi4frag_auto_in_bresp; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_becho_extra_id = axi4frag_auto_in_becho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_arready = axi4frag_auto_in_arready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_rvalid = axi4frag_auto_in_rvalid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_rid = axi4frag_auto_in_rid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_rdata = axi4frag_auto_in_rdata; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_rresp = axi4frag_auto_in_rresp; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_recho_extra_id = axi4frag_auto_in_recho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_rlast = axi4frag_auto_in_rlast; // @[LazyModule.scala 296:16]
  assign axi4yank_1_clock = clock;
  assign axi4yank_1_reset = reset;
  assign axi4yank_1_auto_in_awvalid = axi4index_1_auto_out_awvalid; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_awid = axi4index_1_auto_out_awid; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_awaddr = axi4index_1_auto_out_awaddr; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_awlen = axi4index_1_auto_out_awlen; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_awsize = axi4index_1_auto_out_awsize; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_awburst = axi4index_1_auto_out_awburst; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_awecho_tl_state_size = axi4index_1_auto_out_awecho_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_awecho_tl_state_source = axi4index_1_auto_out_awecho_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_awecho_extra_id = axi4index_1_auto_out_awecho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_wvalid = axi4index_1_auto_out_wvalid; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_wdata = axi4index_1_auto_out_wdata; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_wstrb = axi4index_1_auto_out_wstrb; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_wlast = axi4index_1_auto_out_wlast; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_bready = axi4index_1_auto_out_bready; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_arvalid = axi4index_1_auto_out_arvalid; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_arid = axi4index_1_auto_out_arid; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_araddr = axi4index_1_auto_out_araddr; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_arlen = axi4index_1_auto_out_arlen; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_arsize = axi4index_1_auto_out_arsize; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_arburst = axi4index_1_auto_out_arburst; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_arecho_tl_state_size = axi4index_1_auto_out_arecho_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_arecho_tl_state_source = axi4index_1_auto_out_arecho_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_arecho_extra_id = axi4index_1_auto_out_arecho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_in_rready = axi4index_1_auto_out_rready; // @[LazyModule.scala 296:16]
  assign axi4yank_1_auto_out_awready = master_mem_0_awready; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_wready = master_mem_0_wready; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_bvalid = master_mem_0_bvalid; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_bid = master_mem_0_bid; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_bresp = master_mem_0_bresp; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_arready = master_mem_0_arready; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_rvalid = master_mem_0_rvalid; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_rid = master_mem_0_rid; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_rdata = master_mem_0_rdata; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_rresp = master_mem_0_rresp; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4yank_1_auto_out_rlast = master_mem_0_rlast; // @[Nodes.scala 1210:84 Nodes.scala 1694:56]
  assign axi4index_1_auto_in_awvalid = tl2axi4_auto_out_awvalid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_awid = tl2axi4_auto_out_awid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_awaddr = tl2axi4_auto_out_awaddr; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_awlen = tl2axi4_auto_out_awlen; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_awsize = tl2axi4_auto_out_awsize; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_awburst = tl2axi4_auto_out_awburst; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_awecho_tl_state_size = tl2axi4_auto_out_awecho_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_awecho_tl_state_source = tl2axi4_auto_out_awecho_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_wvalid = tl2axi4_auto_out_wvalid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_wdata = tl2axi4_auto_out_wdata; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_wstrb = tl2axi4_auto_out_wstrb; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_wlast = tl2axi4_auto_out_wlast; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_bready = tl2axi4_auto_out_bready; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_arvalid = tl2axi4_auto_out_arvalid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_arid = tl2axi4_auto_out_arid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_araddr = tl2axi4_auto_out_araddr; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_arlen = tl2axi4_auto_out_arlen; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_arsize = tl2axi4_auto_out_arsize; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_arburst = tl2axi4_auto_out_arburst; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_arecho_tl_state_size = tl2axi4_auto_out_arecho_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_arecho_tl_state_source = tl2axi4_auto_out_arecho_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_in_rready = tl2axi4_auto_out_rready; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_awready = axi4yank_1_auto_in_awready; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_wready = axi4yank_1_auto_in_wready; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_bvalid = axi4yank_1_auto_in_bvalid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_bid = axi4yank_1_auto_in_bid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_bresp = axi4yank_1_auto_in_bresp; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_becho_tl_state_size = axi4yank_1_auto_in_becho_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_becho_tl_state_source = axi4yank_1_auto_in_becho_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_becho_extra_id = axi4yank_1_auto_in_becho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_arready = axi4yank_1_auto_in_arready; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_rvalid = axi4yank_1_auto_in_rvalid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_rid = axi4yank_1_auto_in_rid; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_rdata = axi4yank_1_auto_in_rdata; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_rresp = axi4yank_1_auto_in_rresp; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_recho_tl_state_size = axi4yank_1_auto_in_recho_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_recho_tl_state_source = axi4yank_1_auto_in_recho_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_recho_extra_id = axi4yank_1_auto_in_recho_extra_id; // @[LazyModule.scala 296:16]
  assign axi4index_1_auto_out_rlast = axi4yank_1_auto_in_rlast; // @[LazyModule.scala 296:16]
  assign tl2axi4_clock = clock;
  assign tl2axi4_reset = reset;
  assign tl2axi4_auto_in_a_valid = xbar_auto_out_0_a_valid; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_a_bits_opcode = xbar_auto_out_0_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_a_bits_param = xbar_auto_out_0_a_bits_param; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_a_bits_size = xbar_auto_out_0_a_bits_size; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_a_bits_source = xbar_auto_out_0_a_bits_source; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_a_bits_address = xbar_auto_out_0_a_bits_address; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_a_bits_mask = xbar_auto_out_0_a_bits_mask; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_a_bits_data = xbar_auto_out_0_a_bits_data; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_a_bits_corrupt = xbar_auto_out_0_a_bits_corrupt; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_in_d_ready = xbar_auto_out_0_d_ready; // @[LazyModule.scala 298:16]
  assign tl2axi4_auto_out_awready = axi4index_1_auto_in_awready; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_wready = axi4index_1_auto_in_wready; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_bvalid = axi4index_1_auto_in_bvalid; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_bid = axi4index_1_auto_in_bid; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_bresp = axi4index_1_auto_in_bresp; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_becho_tl_state_size = axi4index_1_auto_in_becho_tl_state_size; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_becho_tl_state_source = axi4index_1_auto_in_becho_tl_state_source; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_arready = axi4index_1_auto_in_arready; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_rvalid = axi4index_1_auto_in_rvalid; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_rid = axi4index_1_auto_in_rid; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_rdata = axi4index_1_auto_in_rdata; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_rresp = axi4index_1_auto_in_rresp; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_recho_tl_state_size = axi4index_1_auto_in_recho_tl_state_size; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_recho_tl_state_source = axi4index_1_auto_in_recho_tl_state_source; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_rlast = axi4index_1_auto_in_rlast; // @[LazyModule.scala 296:16]
  assign err_clock = clock;
  assign err_reset = reset;
  assign err_auto_in_a_valid = widget_2_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign err_auto_in_a_bits_opcode = widget_2_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign err_auto_in_a_bits_param = widget_2_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign err_auto_in_a_bits_size = widget_2_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign err_auto_in_a_bits_source = widget_2_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign err_auto_in_a_bits_address = widget_2_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign err_auto_in_a_bits_mask = widget_2_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign err_auto_in_a_bits_corrupt = widget_2_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16]
  assign err_auto_in_c_valid = widget_2_auto_out_c_valid; // @[LazyModule.scala 296:16]
  assign err_auto_in_c_bits_opcode = widget_2_auto_out_c_bits_opcode; // @[LazyModule.scala 296:16]
  assign err_auto_in_c_bits_param = widget_2_auto_out_c_bits_param; // @[LazyModule.scala 296:16]
  assign err_auto_in_c_bits_size = widget_2_auto_out_c_bits_size; // @[LazyModule.scala 296:16]
  assign err_auto_in_c_bits_source = widget_2_auto_out_c_bits_source; // @[LazyModule.scala 296:16]
  assign err_auto_in_c_bits_address = widget_2_auto_out_c_bits_address; // @[LazyModule.scala 296:16]
  assign err_auto_in_d_ready = widget_2_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign err_auto_in_e_valid = widget_2_auto_out_e_valid; // @[LazyModule.scala 296:16]
  assign atomics_clock = clock;
  assign atomics_reset = reset;
  assign atomics_auto_in_a_valid = fixer_1_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_a_bits_opcode = fixer_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_a_bits_param = fixer_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_a_bits_size = fixer_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_a_bits_source = fixer_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_a_bits_address = fixer_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_a_bits_mask = fixer_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_a_bits_data = fixer_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_c_valid = fixer_1_auto_out_c_valid; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_c_bits_opcode = fixer_1_auto_out_c_bits_opcode; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_c_bits_param = fixer_1_auto_out_c_bits_param; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_c_bits_size = fixer_1_auto_out_c_bits_size; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_c_bits_source = fixer_1_auto_out_c_bits_source; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_c_bits_address = fixer_1_auto_out_c_bits_address; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_d_ready = fixer_1_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_e_valid = fixer_1_auto_out_e_valid; // @[LazyModule.scala 296:16]
  assign atomics_auto_in_e_bits_sink = fixer_1_auto_out_e_bits_sink; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_a_ready = xbar_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_c_ready = xbar_auto_in_c_ready; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_valid = xbar_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_opcode = xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_param = xbar_auto_in_d_bits_param; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_size = xbar_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_source = xbar_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_denied = xbar_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_data = xbar_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_corrupt = xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_e_ready = xbar_auto_in_e_ready; // @[LazyModule.scala 296:16]
  assign fixer_1_clock = clock;
  assign fixer_1_reset = reset;
  assign fixer_1_auto_in_a_valid = hints_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_a_bits_opcode = hints_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_a_bits_param = hints_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_a_bits_size = hints_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_a_bits_source = hints_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_a_bits_address = hints_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_a_bits_mask = hints_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_a_bits_data = hints_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_c_valid = hints_auto_out_c_valid; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_c_bits_opcode = hints_auto_out_c_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_c_bits_param = hints_auto_out_c_bits_param; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_c_bits_size = hints_auto_out_c_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_c_bits_source = hints_auto_out_c_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_c_bits_address = hints_auto_out_c_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_d_ready = hints_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_e_valid = hints_auto_out_e_valid; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_in_e_bits_sink = hints_auto_out_e_bits_sink; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_a_ready = atomics_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_c_ready = atomics_auto_in_c_ready; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_d_valid = atomics_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_d_bits_opcode = atomics_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_d_bits_param = atomics_auto_in_d_bits_param; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_d_bits_size = atomics_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_d_bits_source = atomics_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_d_bits_denied = atomics_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_d_bits_data = atomics_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_d_bits_corrupt = atomics_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign fixer_1_auto_out_e_ready = atomics_auto_in_e_ready; // @[LazyModule.scala 296:16]
  assign hints_clock = clock;
  assign hints_reset = reset;
  assign hints_auto_in_a_valid = widget_1_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign hints_auto_in_a_bits_opcode = widget_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign hints_auto_in_a_bits_param = widget_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign hints_auto_in_a_bits_size = widget_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign hints_auto_in_a_bits_source = widget_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign hints_auto_in_a_bits_address = widget_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign hints_auto_in_a_bits_mask = widget_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign hints_auto_in_a_bits_data = widget_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign hints_auto_in_c_valid = widget_1_auto_out_c_valid; // @[LazyModule.scala 296:16]
  assign hints_auto_in_c_bits_opcode = widget_1_auto_out_c_bits_opcode; // @[LazyModule.scala 296:16]
  assign hints_auto_in_c_bits_param = widget_1_auto_out_c_bits_param; // @[LazyModule.scala 296:16]
  assign hints_auto_in_c_bits_size = widget_1_auto_out_c_bits_size; // @[LazyModule.scala 296:16]
  assign hints_auto_in_c_bits_source = widget_1_auto_out_c_bits_source; // @[LazyModule.scala 296:16]
  assign hints_auto_in_c_bits_address = widget_1_auto_out_c_bits_address; // @[LazyModule.scala 296:16]
  assign hints_auto_in_d_ready = widget_1_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign hints_auto_in_e_valid = widget_1_auto_out_e_valid; // @[LazyModule.scala 296:16]
  assign hints_auto_in_e_bits_sink = widget_1_auto_out_e_bits_sink; // @[LazyModule.scala 296:16]
  assign hints_auto_out_a_ready = fixer_1_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign hints_auto_out_c_ready = fixer_1_auto_in_c_ready; // @[LazyModule.scala 296:16]
  assign hints_auto_out_d_valid = fixer_1_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign hints_auto_out_d_bits_opcode = fixer_1_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign hints_auto_out_d_bits_param = fixer_1_auto_in_d_bits_param; // @[LazyModule.scala 296:16]
  assign hints_auto_out_d_bits_size = fixer_1_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign hints_auto_out_d_bits_source = fixer_1_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign hints_auto_out_d_bits_denied = fixer_1_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign hints_auto_out_d_bits_data = fixer_1_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign hints_auto_out_d_bits_corrupt = fixer_1_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign hints_auto_out_e_ready = fixer_1_auto_in_e_ready; // @[LazyModule.scala 296:16]
  assign widget_1_clock = clock;
  assign widget_1_reset = reset;
  assign widget_1_auto_in_a_valid = chiplink_auto_mbypass_out_a_valid; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_a_bits_opcode = chiplink_auto_mbypass_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_a_bits_param = chiplink_auto_mbypass_out_a_bits_param; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_a_bits_size = chiplink_auto_mbypass_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_a_bits_source = chiplink_auto_mbypass_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_a_bits_address = chiplink_auto_mbypass_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_a_bits_mask = chiplink_auto_mbypass_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_a_bits_data = chiplink_auto_mbypass_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_c_valid = chiplink_auto_mbypass_out_c_valid; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_c_bits_opcode = chiplink_auto_mbypass_out_c_bits_opcode; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_c_bits_param = chiplink_auto_mbypass_out_c_bits_param; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_c_bits_size = chiplink_auto_mbypass_out_c_bits_size; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_c_bits_source = chiplink_auto_mbypass_out_c_bits_source; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_c_bits_address = chiplink_auto_mbypass_out_c_bits_address; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_d_ready = chiplink_auto_mbypass_out_d_ready; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_e_valid = chiplink_auto_mbypass_out_e_valid; // @[LazyModule.scala 298:16]
  assign widget_1_auto_in_e_bits_sink = chiplink_auto_mbypass_out_e_bits_sink; // @[LazyModule.scala 298:16]
  assign widget_1_auto_out_a_ready = hints_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_c_ready = hints_auto_in_c_ready; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_d_valid = hints_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_d_bits_opcode = hints_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_d_bits_param = hints_auto_in_d_bits_param; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_d_bits_size = hints_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_d_bits_source = hints_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_d_bits_denied = hints_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_d_bits_data = hints_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_d_bits_corrupt = hints_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign widget_1_auto_out_e_ready = hints_auto_in_e_ready; // @[LazyModule.scala 296:16]
  assign widget_2_clock = clock;
  assign widget_2_reset = reset;
  assign widget_2_auto_in_a_valid = xbar_auto_out_1_a_valid; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_a_bits_opcode = xbar_auto_out_1_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_a_bits_param = xbar_auto_out_1_a_bits_param; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_a_bits_size = xbar_auto_out_1_a_bits_size; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_a_bits_source = xbar_auto_out_1_a_bits_source; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_a_bits_address = xbar_auto_out_1_a_bits_address; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_a_bits_mask = xbar_auto_out_1_a_bits_mask; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_a_bits_corrupt = xbar_auto_out_1_a_bits_corrupt; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_c_valid = xbar_auto_out_1_c_valid; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_c_bits_opcode = xbar_auto_out_1_c_bits_opcode; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_c_bits_param = xbar_auto_out_1_c_bits_param; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_c_bits_size = xbar_auto_out_1_c_bits_size; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_c_bits_source = xbar_auto_out_1_c_bits_source; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_c_bits_address = xbar_auto_out_1_c_bits_address; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_d_ready = xbar_auto_out_1_d_ready; // @[LazyModule.scala 298:16]
  assign widget_2_auto_in_e_valid = xbar_auto_out_1_e_valid; // @[LazyModule.scala 298:16]
  assign widget_2_auto_out_a_ready = err_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign widget_2_auto_out_c_ready = err_auto_in_c_ready; // @[LazyModule.scala 296:16]
  assign widget_2_auto_out_d_valid = err_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign widget_2_auto_out_d_bits_opcode = err_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_2_auto_out_d_bits_param = err_auto_in_d_bits_param; // @[LazyModule.scala 296:16]
  assign widget_2_auto_out_d_bits_size = err_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign widget_2_auto_out_d_bits_source = err_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign widget_2_auto_out_d_bits_denied = err_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign widget_2_auto_out_d_bits_corrupt = err_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
endmodule
module ChipLinkBridgeLazy(
  input         clock,
  input         reset,
  input         io_master_awready,
  output        io_master_awvalid,
  output [3:0]  io_master_awid,
  output [31:0] io_master_awaddr,
  output [7:0]  io_master_awlen,
  output [2:0]  io_master_awsize,
  output [1:0]  io_master_awburst,
  input         io_master_wready,
  output        io_master_wvalid,
  output [63:0] io_master_wdata,
  output [7:0]  io_master_wstrb,
  output        io_master_wlast,
  output        io_master_bready,
  input         io_master_bvalid,
  input  [3:0]  io_master_bid,
  input  [1:0]  io_master_bresp,
  input         io_master_arready,
  output        io_master_arvalid,
  output [3:0]  io_master_arid,
  output [31:0] io_master_araddr,
  output [7:0]  io_master_arlen,
  output [2:0]  io_master_arsize,
  output [1:0]  io_master_arburst,
  output        io_master_rready,
  input         io_master_rvalid,
  input  [3:0]  io_master_rid,
  input  [63:0] io_master_rdata,
  input  [1:0]  io_master_rresp,
  input         io_master_rlast,
  output        io_slave_awready,
  input         io_slave_awvalid,
  input  [3:0]  io_slave_awid,
  input  [31:0] io_slave_awaddr,
  input  [7:0]  io_slave_awlen,
  input  [2:0]  io_slave_awsize,
  input  [1:0]  io_slave_awburst,
  output        io_slave_wready,
  input         io_slave_wvalid,
  input  [63:0] io_slave_wdata,
  input  [7:0]  io_slave_wstrb,
  input         io_slave_wlast,
  input         io_slave_bready,
  output        io_slave_bvalid,
  output [3:0]  io_slave_bid,
  output [1:0]  io_slave_bresp,
  output        io_slave_arready,
  input         io_slave_arvalid,
  input  [3:0]  io_slave_arid,
  input  [31:0] io_slave_araddr,
  input  [7:0]  io_slave_arlen,
  input  [2:0]  io_slave_arsize,
  input  [1:0]  io_slave_arburst,
  input         io_slave_rready,
  output        io_slave_rvalid,
  output [3:0]  io_slave_rid,
  output [63:0] io_slave_rdata,
  output [1:0]  io_slave_rresp,
  output        io_slave_rlast,
  output        fpga_io_c2b_clk,
  output        fpga_io_c2b_rst,
  output        fpga_io_c2b_send,
  output [7:0]  fpga_io_c2b_data,
  input         fpga_io_b2c_clk,
  input         fpga_io_b2c_rst,
  input         fpga_io_b2c_send,
  input  [7:0]  fpga_io_b2c_data
);
  wire  chipLinkConverter_clock; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_reset; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_awready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_awvalid; // @[TestHarness.scala 44:37]
  wire [3:0] chipLinkConverter_slave_0_awid; // @[TestHarness.scala 44:37]
  wire [31:0] chipLinkConverter_slave_0_awaddr; // @[TestHarness.scala 44:37]
  wire [7:0] chipLinkConverter_slave_0_awlen; // @[TestHarness.scala 44:37]
  wire [2:0] chipLinkConverter_slave_0_awsize; // @[TestHarness.scala 44:37]
  wire [1:0] chipLinkConverter_slave_0_awburst; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_wready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_wvalid; // @[TestHarness.scala 44:37]
  wire [63:0] chipLinkConverter_slave_0_wdata; // @[TestHarness.scala 44:37]
  wire [7:0] chipLinkConverter_slave_0_wstrb; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_wlast; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_bready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_bvalid; // @[TestHarness.scala 44:37]
  wire [3:0] chipLinkConverter_slave_0_bid; // @[TestHarness.scala 44:37]
  wire [1:0] chipLinkConverter_slave_0_bresp; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_arready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_arvalid; // @[TestHarness.scala 44:37]
  wire [3:0] chipLinkConverter_slave_0_arid; // @[TestHarness.scala 44:37]
  wire [31:0] chipLinkConverter_slave_0_araddr; // @[TestHarness.scala 44:37]
  wire [7:0] chipLinkConverter_slave_0_arlen; // @[TestHarness.scala 44:37]
  wire [2:0] chipLinkConverter_slave_0_arsize; // @[TestHarness.scala 44:37]
  wire [1:0] chipLinkConverter_slave_0_arburst; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_rready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_rvalid; // @[TestHarness.scala 44:37]
  wire [3:0] chipLinkConverter_slave_0_rid; // @[TestHarness.scala 44:37]
  wire [63:0] chipLinkConverter_slave_0_rdata; // @[TestHarness.scala 44:37]
  wire [1:0] chipLinkConverter_slave_0_rresp; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_slave_0_rlast; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_awready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_awvalid; // @[TestHarness.scala 44:37]
  wire [3:0] chipLinkConverter_master_mem_0_awid; // @[TestHarness.scala 44:37]
  wire [31:0] chipLinkConverter_master_mem_0_awaddr; // @[TestHarness.scala 44:37]
  wire [7:0] chipLinkConverter_master_mem_0_awlen; // @[TestHarness.scala 44:37]
  wire [2:0] chipLinkConverter_master_mem_0_awsize; // @[TestHarness.scala 44:37]
  wire [1:0] chipLinkConverter_master_mem_0_awburst; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_wready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_wvalid; // @[TestHarness.scala 44:37]
  wire [63:0] chipLinkConverter_master_mem_0_wdata; // @[TestHarness.scala 44:37]
  wire [7:0] chipLinkConverter_master_mem_0_wstrb; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_wlast; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_bready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_bvalid; // @[TestHarness.scala 44:37]
  wire [3:0] chipLinkConverter_master_mem_0_bid; // @[TestHarness.scala 44:37]
  wire [1:0] chipLinkConverter_master_mem_0_bresp; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_arready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_arvalid; // @[TestHarness.scala 44:37]
  wire [3:0] chipLinkConverter_master_mem_0_arid; // @[TestHarness.scala 44:37]
  wire [31:0] chipLinkConverter_master_mem_0_araddr; // @[TestHarness.scala 44:37]
  wire [7:0] chipLinkConverter_master_mem_0_arlen; // @[TestHarness.scala 44:37]
  wire [2:0] chipLinkConverter_master_mem_0_arsize; // @[TestHarness.scala 44:37]
  wire [1:0] chipLinkConverter_master_mem_0_arburst; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_rready; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_rvalid; // @[TestHarness.scala 44:37]
  wire [3:0] chipLinkConverter_master_mem_0_rid; // @[TestHarness.scala 44:37]
  wire [63:0] chipLinkConverter_master_mem_0_rdata; // @[TestHarness.scala 44:37]
  wire [1:0] chipLinkConverter_master_mem_0_rresp; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_master_mem_0_rlast; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_fpga_io_c2b_clk; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_fpga_io_c2b_rst; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_fpga_io_c2b_send; // @[TestHarness.scala 44:37]
  wire [7:0] chipLinkConverter_fpga_io_c2b_data; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_fpga_io_b2c_clk; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_fpga_io_b2c_rst; // @[TestHarness.scala 44:37]
  wire  chipLinkConverter_fpga_io_b2c_send; // @[TestHarness.scala 44:37]
  wire [7:0] chipLinkConverter_fpga_io_b2c_data; // @[TestHarness.scala 44:37]
  ChipLinkMaster chipLinkConverter ( // @[TestHarness.scala 44:37]
    .clock(chipLinkConverter_clock),
    .reset(chipLinkConverter_reset),
    .slave_0_awready(chipLinkConverter_slave_0_awready),
    .slave_0_awvalid(chipLinkConverter_slave_0_awvalid),
    .slave_0_awid(chipLinkConverter_slave_0_awid),
    .slave_0_awaddr(chipLinkConverter_slave_0_awaddr),
    .slave_0_awlen(chipLinkConverter_slave_0_awlen),
    .slave_0_awsize(chipLinkConverter_slave_0_awsize),
    .slave_0_awburst(chipLinkConverter_slave_0_awburst),
    .slave_0_wready(chipLinkConverter_slave_0_wready),
    .slave_0_wvalid(chipLinkConverter_slave_0_wvalid),
    .slave_0_wdata(chipLinkConverter_slave_0_wdata),
    .slave_0_wstrb(chipLinkConverter_slave_0_wstrb),
    .slave_0_wlast(chipLinkConverter_slave_0_wlast),
    .slave_0_bready(chipLinkConverter_slave_0_bready),
    .slave_0_bvalid(chipLinkConverter_slave_0_bvalid),
    .slave_0_bid(chipLinkConverter_slave_0_bid),
    .slave_0_bresp(chipLinkConverter_slave_0_bresp),
    .slave_0_arready(chipLinkConverter_slave_0_arready),
    .slave_0_arvalid(chipLinkConverter_slave_0_arvalid),
    .slave_0_arid(chipLinkConverter_slave_0_arid),
    .slave_0_araddr(chipLinkConverter_slave_0_araddr),
    .slave_0_arlen(chipLinkConverter_slave_0_arlen),
    .slave_0_arsize(chipLinkConverter_slave_0_arsize),
    .slave_0_arburst(chipLinkConverter_slave_0_arburst),
    .slave_0_rready(chipLinkConverter_slave_0_rready),
    .slave_0_rvalid(chipLinkConverter_slave_0_rvalid),
    .slave_0_rid(chipLinkConverter_slave_0_rid),
    .slave_0_rdata(chipLinkConverter_slave_0_rdata),
    .slave_0_rresp(chipLinkConverter_slave_0_rresp),
    .slave_0_rlast(chipLinkConverter_slave_0_rlast),
    .master_mem_0_awready(chipLinkConverter_master_mem_0_awready),
    .master_mem_0_awvalid(chipLinkConverter_master_mem_0_awvalid),
    .master_mem_0_awid(chipLinkConverter_master_mem_0_awid),
    .master_mem_0_awaddr(chipLinkConverter_master_mem_0_awaddr),
    .master_mem_0_awlen(chipLinkConverter_master_mem_0_awlen),
    .master_mem_0_awsize(chipLinkConverter_master_mem_0_awsize),
    .master_mem_0_awburst(chipLinkConverter_master_mem_0_awburst),
    .master_mem_0_wready(chipLinkConverter_master_mem_0_wready),
    .master_mem_0_wvalid(chipLinkConverter_master_mem_0_wvalid),
    .master_mem_0_wdata(chipLinkConverter_master_mem_0_wdata),
    .master_mem_0_wstrb(chipLinkConverter_master_mem_0_wstrb),
    .master_mem_0_wlast(chipLinkConverter_master_mem_0_wlast),
    .master_mem_0_bready(chipLinkConverter_master_mem_0_bready),
    .master_mem_0_bvalid(chipLinkConverter_master_mem_0_bvalid),
    .master_mem_0_bid(chipLinkConverter_master_mem_0_bid),
    .master_mem_0_bresp(chipLinkConverter_master_mem_0_bresp),
    .master_mem_0_arready(chipLinkConverter_master_mem_0_arready),
    .master_mem_0_arvalid(chipLinkConverter_master_mem_0_arvalid),
    .master_mem_0_arid(chipLinkConverter_master_mem_0_arid),
    .master_mem_0_araddr(chipLinkConverter_master_mem_0_araddr),
    .master_mem_0_arlen(chipLinkConverter_master_mem_0_arlen),
    .master_mem_0_arsize(chipLinkConverter_master_mem_0_arsize),
    .master_mem_0_arburst(chipLinkConverter_master_mem_0_arburst),
    .master_mem_0_rready(chipLinkConverter_master_mem_0_rready),
    .master_mem_0_rvalid(chipLinkConverter_master_mem_0_rvalid),
    .master_mem_0_rid(chipLinkConverter_master_mem_0_rid),
    .master_mem_0_rdata(chipLinkConverter_master_mem_0_rdata),
    .master_mem_0_rresp(chipLinkConverter_master_mem_0_rresp),
    .master_mem_0_rlast(chipLinkConverter_master_mem_0_rlast),
    .fpga_io_c2b_clk(chipLinkConverter_fpga_io_c2b_clk),
    .fpga_io_c2b_rst(chipLinkConverter_fpga_io_c2b_rst),
    .fpga_io_c2b_send(chipLinkConverter_fpga_io_c2b_send),
    .fpga_io_c2b_data(chipLinkConverter_fpga_io_c2b_data),
    .fpga_io_b2c_clk(chipLinkConverter_fpga_io_b2c_clk),
    .fpga_io_b2c_rst(chipLinkConverter_fpga_io_b2c_rst),
    .fpga_io_b2c_send(chipLinkConverter_fpga_io_b2c_send),
    .fpga_io_b2c_data(chipLinkConverter_fpga_io_b2c_data)
  );
  assign io_master_awvalid = chipLinkConverter_master_mem_0_awvalid; // @[TestHarness.scala 51:15]
  assign io_master_awid = chipLinkConverter_master_mem_0_awid; // @[TestHarness.scala 51:15]
  assign io_master_awaddr = chipLinkConverter_master_mem_0_awaddr; // @[TestHarness.scala 51:15]
  assign io_master_awlen = chipLinkConverter_master_mem_0_awlen; // @[TestHarness.scala 51:15]
  assign io_master_awsize = chipLinkConverter_master_mem_0_awsize; // @[TestHarness.scala 51:15]
  assign io_master_awburst = chipLinkConverter_master_mem_0_awburst; // @[TestHarness.scala 51:15]
  assign io_master_wvalid = chipLinkConverter_master_mem_0_wvalid; // @[TestHarness.scala 51:15]
  assign io_master_wdata = chipLinkConverter_master_mem_0_wdata; // @[TestHarness.scala 51:15]
  assign io_master_wstrb = chipLinkConverter_master_mem_0_wstrb; // @[TestHarness.scala 51:15]
  assign io_master_wlast = chipLinkConverter_master_mem_0_wlast; // @[TestHarness.scala 51:15]
  assign io_master_bready = chipLinkConverter_master_mem_0_bready; // @[TestHarness.scala 51:15]
  assign io_master_arvalid = chipLinkConverter_master_mem_0_arvalid; // @[TestHarness.scala 51:15]
  assign io_master_arid = chipLinkConverter_master_mem_0_arid; // @[TestHarness.scala 51:15]
  assign io_master_araddr = chipLinkConverter_master_mem_0_araddr; // @[TestHarness.scala 51:15]
  assign io_master_arlen = chipLinkConverter_master_mem_0_arlen; // @[TestHarness.scala 51:15]
  assign io_master_arsize = chipLinkConverter_master_mem_0_arsize; // @[TestHarness.scala 51:15]
  assign io_master_arburst = chipLinkConverter_master_mem_0_arburst; // @[TestHarness.scala 51:15]
  assign io_master_rready = chipLinkConverter_master_mem_0_rready; // @[TestHarness.scala 51:15]
  assign io_slave_awready = chipLinkConverter_slave_0_awready; // @[TestHarness.scala 50:34]
  assign io_slave_wready = chipLinkConverter_slave_0_wready; // @[TestHarness.scala 50:34]
  assign io_slave_bvalid = chipLinkConverter_slave_0_bvalid; // @[TestHarness.scala 50:34]
  assign io_slave_bid = chipLinkConverter_slave_0_bid; // @[TestHarness.scala 50:34]
  assign io_slave_bresp = chipLinkConverter_slave_0_bresp; // @[TestHarness.scala 50:34]
  assign io_slave_arready = chipLinkConverter_slave_0_arready; // @[TestHarness.scala 50:34]
  assign io_slave_rvalid = chipLinkConverter_slave_0_rvalid; // @[TestHarness.scala 50:34]
  assign io_slave_rid = chipLinkConverter_slave_0_rid; // @[TestHarness.scala 50:34]
  assign io_slave_rdata = chipLinkConverter_slave_0_rdata; // @[TestHarness.scala 50:34]
  assign io_slave_rresp = chipLinkConverter_slave_0_rresp; // @[TestHarness.scala 50:34]
  assign io_slave_rlast = chipLinkConverter_slave_0_rlast; // @[TestHarness.scala 50:34]
  assign fpga_io_c2b_clk = chipLinkConverter_fpga_io_c2b_clk; // @[TestHarness.scala 49:13]
  assign fpga_io_c2b_rst = chipLinkConverter_fpga_io_c2b_rst; // @[TestHarness.scala 49:13]
  assign fpga_io_c2b_send = chipLinkConverter_fpga_io_c2b_send; // @[TestHarness.scala 49:13]
  assign fpga_io_c2b_data = chipLinkConverter_fpga_io_c2b_data; // @[TestHarness.scala 49:13]
  assign chipLinkConverter_clock = clock;
  assign chipLinkConverter_reset = reset;
  assign chipLinkConverter_slave_0_awvalid = io_slave_awvalid; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_awid = io_slave_awid; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_awaddr = io_slave_awaddr; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_awlen = io_slave_awlen; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_awsize = io_slave_awsize; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_awburst = io_slave_awburst; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_wvalid = io_slave_wvalid; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_wdata = io_slave_wdata; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_wstrb = io_slave_wstrb; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_wlast = io_slave_wlast; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_bready = io_slave_bready; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_arvalid = io_slave_arvalid; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_arid = io_slave_arid; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_araddr = io_slave_araddr; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_arlen = io_slave_arlen; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_arsize = io_slave_arsize; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_arburst = io_slave_arburst; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_slave_0_rready = io_slave_rready; // @[TestHarness.scala 50:34]
  assign chipLinkConverter_master_mem_0_awready = io_master_awready; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_wready = io_master_wready; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_bvalid = io_master_bvalid; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_bid = io_master_bid; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_bresp = io_master_bresp; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_arready = io_master_arready; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_rvalid = io_master_rvalid; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_rid = io_master_rid; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_rdata = io_master_rdata; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_rresp = io_master_rresp; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_master_mem_0_rlast = io_master_rlast; // @[TestHarness.scala 51:15]
  assign chipLinkConverter_fpga_io_b2c_clk = fpga_io_b2c_clk; // @[TestHarness.scala 49:13]
  assign chipLinkConverter_fpga_io_b2c_rst = fpga_io_b2c_rst; // @[TestHarness.scala 49:13]
  assign chipLinkConverter_fpga_io_b2c_send = fpga_io_b2c_send; // @[TestHarness.scala 49:13]
  assign chipLinkConverter_fpga_io_b2c_data = fpga_io_b2c_data; // @[TestHarness.scala 49:13]
endmodule
module ChiplinkBridge(
  input         clock,
  input         reset,
  input         mem_axi4_0_awready,
  output        mem_axi4_0_awvalid,
  output [3:0]  mem_axi4_0_awid,
  output [31:0] mem_axi4_0_awaddr,
  output [7:0]  mem_axi4_0_awlen,
  output [2:0]  mem_axi4_0_awsize,
  output [1:0]  mem_axi4_0_awburst,
  input         mem_axi4_0_wready,
  output        mem_axi4_0_wvalid,
  output [63:0] mem_axi4_0_wdata,
  output [7:0]  mem_axi4_0_wstrb,
  output        mem_axi4_0_wlast,
  output        mem_axi4_0_bready,
  input         mem_axi4_0_bvalid,
  input  [3:0]  mem_axi4_0_bid,
  input  [1:0]  mem_axi4_0_bresp,
  input         mem_axi4_0_arready,
  output        mem_axi4_0_arvalid,
  output [3:0]  mem_axi4_0_arid,
  output [31:0] mem_axi4_0_araddr,
  output [7:0]  mem_axi4_0_arlen,
  output [2:0]  mem_axi4_0_arsize,
  output [1:0]  mem_axi4_0_arburst,
  output        mem_axi4_0_rready,
  input         mem_axi4_0_rvalid,
  input  [3:0]  mem_axi4_0_rid,
  input  [63:0] mem_axi4_0_rdata,
  input  [1:0]  mem_axi4_0_rresp,
  input         mem_axi4_0_rlast,
  output        slave_axi4_mem_0_awready,
  input         slave_axi4_mem_0_awvalid,
  input  [3:0]  slave_axi4_mem_0_awid,
  input  [31:0] slave_axi4_mem_0_awaddr,
  input  [7:0]  slave_axi4_mem_0_awlen,
  input  [2:0]  slave_axi4_mem_0_awsize,
  input  [1:0]  slave_axi4_mem_0_awburst,
  output        slave_axi4_mem_0_wready,
  input         slave_axi4_mem_0_wvalid,
  input  [63:0] slave_axi4_mem_0_wdata,
  input  [7:0]  slave_axi4_mem_0_wstrb,
  input         slave_axi4_mem_0_wlast,
  input         slave_axi4_mem_0_bready,
  output        slave_axi4_mem_0_bvalid,
  output [3:0]  slave_axi4_mem_0_bid,
  output [1:0]  slave_axi4_mem_0_bresp,
  output        slave_axi4_mem_0_arready,
  input         slave_axi4_mem_0_arvalid,
  input  [3:0]  slave_axi4_mem_0_arid,
  input  [31:0] slave_axi4_mem_0_araddr,
  input  [7:0]  slave_axi4_mem_0_arlen,
  input  [2:0]  slave_axi4_mem_0_arsize,
  input  [1:0]  slave_axi4_mem_0_arburst,
  input         slave_axi4_mem_0_rready,
  output        slave_axi4_mem_0_rvalid,
  output [3:0]  slave_axi4_mem_0_rid,
  output [63:0] slave_axi4_mem_0_rdata,
  output [1:0]  slave_axi4_mem_0_rresp,
  output        slave_axi4_mem_0_rlast,
  output        fpga_io_c2b_clk,
  output        fpga_io_c2b_rst,
  output        fpga_io_c2b_send,
  output [7:0]  fpga_io_c2b_data,
  input         fpga_io_b2c_clk,
  input         fpga_io_b2c_rst,
  input         fpga_io_b2c_send,
  input  [7:0]  fpga_io_b2c_data
);
  wire  clBridge_clock; // @[TestHarness.scala 37:25]
  wire  clBridge_reset; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_awready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_awvalid; // @[TestHarness.scala 37:25]
  wire [3:0] clBridge_io_master_awid; // @[TestHarness.scala 37:25]
  wire [31:0] clBridge_io_master_awaddr; // @[TestHarness.scala 37:25]
  wire [7:0] clBridge_io_master_awlen; // @[TestHarness.scala 37:25]
  wire [2:0] clBridge_io_master_awsize; // @[TestHarness.scala 37:25]
  wire [1:0] clBridge_io_master_awburst; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_wready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_wvalid; // @[TestHarness.scala 37:25]
  wire [63:0] clBridge_io_master_wdata; // @[TestHarness.scala 37:25]
  wire [7:0] clBridge_io_master_wstrb; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_wlast; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_bready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_bvalid; // @[TestHarness.scala 37:25]
  wire [3:0] clBridge_io_master_bid; // @[TestHarness.scala 37:25]
  wire [1:0] clBridge_io_master_bresp; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_arready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_arvalid; // @[TestHarness.scala 37:25]
  wire [3:0] clBridge_io_master_arid; // @[TestHarness.scala 37:25]
  wire [31:0] clBridge_io_master_araddr; // @[TestHarness.scala 37:25]
  wire [7:0] clBridge_io_master_arlen; // @[TestHarness.scala 37:25]
  wire [2:0] clBridge_io_master_arsize; // @[TestHarness.scala 37:25]
  wire [1:0] clBridge_io_master_arburst; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_rready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_rvalid; // @[TestHarness.scala 37:25]
  wire [3:0] clBridge_io_master_rid; // @[TestHarness.scala 37:25]
  wire [63:0] clBridge_io_master_rdata; // @[TestHarness.scala 37:25]
  wire [1:0] clBridge_io_master_rresp; // @[TestHarness.scala 37:25]
  wire  clBridge_io_master_rlast; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_awready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_awvalid; // @[TestHarness.scala 37:25]
  wire [3:0] clBridge_io_slave_awid; // @[TestHarness.scala 37:25]
  wire [31:0] clBridge_io_slave_awaddr; // @[TestHarness.scala 37:25]
  wire [7:0] clBridge_io_slave_awlen; // @[TestHarness.scala 37:25]
  wire [2:0] clBridge_io_slave_awsize; // @[TestHarness.scala 37:25]
  wire [1:0] clBridge_io_slave_awburst; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_wready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_wvalid; // @[TestHarness.scala 37:25]
  wire [63:0] clBridge_io_slave_wdata; // @[TestHarness.scala 37:25]
  wire [7:0] clBridge_io_slave_wstrb; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_wlast; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_bready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_bvalid; // @[TestHarness.scala 37:25]
  wire [3:0] clBridge_io_slave_bid; // @[TestHarness.scala 37:25]
  wire [1:0] clBridge_io_slave_bresp; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_arready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_arvalid; // @[TestHarness.scala 37:25]
  wire [3:0] clBridge_io_slave_arid; // @[TestHarness.scala 37:25]
  wire [31:0] clBridge_io_slave_araddr; // @[TestHarness.scala 37:25]
  wire [7:0] clBridge_io_slave_arlen; // @[TestHarness.scala 37:25]
  wire [2:0] clBridge_io_slave_arsize; // @[TestHarness.scala 37:25]
  wire [1:0] clBridge_io_slave_arburst; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_rready; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_rvalid; // @[TestHarness.scala 37:25]
  wire [3:0] clBridge_io_slave_rid; // @[TestHarness.scala 37:25]
  wire [63:0] clBridge_io_slave_rdata; // @[TestHarness.scala 37:25]
  wire [1:0] clBridge_io_slave_rresp; // @[TestHarness.scala 37:25]
  wire  clBridge_io_slave_rlast; // @[TestHarness.scala 37:25]
  wire  clBridge_fpga_io_c2b_clk; // @[TestHarness.scala 37:25]
  wire  clBridge_fpga_io_c2b_rst; // @[TestHarness.scala 37:25]
  wire  clBridge_fpga_io_c2b_send; // @[TestHarness.scala 37:25]
  wire [7:0] clBridge_fpga_io_c2b_data; // @[TestHarness.scala 37:25]
  wire  clBridge_fpga_io_b2c_clk; // @[TestHarness.scala 37:25]
  wire  clBridge_fpga_io_b2c_rst; // @[TestHarness.scala 37:25]
  wire  clBridge_fpga_io_b2c_send; // @[TestHarness.scala 37:25]
  wire [7:0] clBridge_fpga_io_b2c_data; // @[TestHarness.scala 37:25]
  ChipLinkBridgeLazy clBridge ( // @[TestHarness.scala 37:25]
    .clock(clBridge_clock),
    .reset(clBridge_reset),
    .io_master_awready(clBridge_io_master_awready),
    .io_master_awvalid(clBridge_io_master_awvalid),
    .io_master_awid(clBridge_io_master_awid),
    .io_master_awaddr(clBridge_io_master_awaddr),
    .io_master_awlen(clBridge_io_master_awlen),
    .io_master_awsize(clBridge_io_master_awsize),
    .io_master_awburst(clBridge_io_master_awburst),
    .io_master_wready(clBridge_io_master_wready),
    .io_master_wvalid(clBridge_io_master_wvalid),
    .io_master_wdata(clBridge_io_master_wdata),
    .io_master_wstrb(clBridge_io_master_wstrb),
    .io_master_wlast(clBridge_io_master_wlast),
    .io_master_bready(clBridge_io_master_bready),
    .io_master_bvalid(clBridge_io_master_bvalid),
    .io_master_bid(clBridge_io_master_bid),
    .io_master_bresp(clBridge_io_master_bresp),
    .io_master_arready(clBridge_io_master_arready),
    .io_master_arvalid(clBridge_io_master_arvalid),
    .io_master_arid(clBridge_io_master_arid),
    .io_master_araddr(clBridge_io_master_araddr),
    .io_master_arlen(clBridge_io_master_arlen),
    .io_master_arsize(clBridge_io_master_arsize),
    .io_master_arburst(clBridge_io_master_arburst),
    .io_master_rready(clBridge_io_master_rready),
    .io_master_rvalid(clBridge_io_master_rvalid),
    .io_master_rid(clBridge_io_master_rid),
    .io_master_rdata(clBridge_io_master_rdata),
    .io_master_rresp(clBridge_io_master_rresp),
    .io_master_rlast(clBridge_io_master_rlast),
    .io_slave_awready(clBridge_io_slave_awready),
    .io_slave_awvalid(clBridge_io_slave_awvalid),
    .io_slave_awid(clBridge_io_slave_awid),
    .io_slave_awaddr(clBridge_io_slave_awaddr),
    .io_slave_awlen(clBridge_io_slave_awlen),
    .io_slave_awsize(clBridge_io_slave_awsize),
    .io_slave_awburst(clBridge_io_slave_awburst),
    .io_slave_wready(clBridge_io_slave_wready),
    .io_slave_wvalid(clBridge_io_slave_wvalid),
    .io_slave_wdata(clBridge_io_slave_wdata),
    .io_slave_wstrb(clBridge_io_slave_wstrb),
    .io_slave_wlast(clBridge_io_slave_wlast),
    .io_slave_bready(clBridge_io_slave_bready),
    .io_slave_bvalid(clBridge_io_slave_bvalid),
    .io_slave_bid(clBridge_io_slave_bid),
    .io_slave_bresp(clBridge_io_slave_bresp),
    .io_slave_arready(clBridge_io_slave_arready),
    .io_slave_arvalid(clBridge_io_slave_arvalid),
    .io_slave_arid(clBridge_io_slave_arid),
    .io_slave_araddr(clBridge_io_slave_araddr),
    .io_slave_arlen(clBridge_io_slave_arlen),
    .io_slave_arsize(clBridge_io_slave_arsize),
    .io_slave_arburst(clBridge_io_slave_arburst),
    .io_slave_rready(clBridge_io_slave_rready),
    .io_slave_rvalid(clBridge_io_slave_rvalid),
    .io_slave_rid(clBridge_io_slave_rid),
    .io_slave_rdata(clBridge_io_slave_rdata),
    .io_slave_rresp(clBridge_io_slave_rresp),
    .io_slave_rlast(clBridge_io_slave_rlast),
    .fpga_io_c2b_clk(clBridge_fpga_io_c2b_clk),
    .fpga_io_c2b_rst(clBridge_fpga_io_c2b_rst),
    .fpga_io_c2b_send(clBridge_fpga_io_c2b_send),
    .fpga_io_c2b_data(clBridge_fpga_io_c2b_data),
    .fpga_io_b2c_clk(clBridge_fpga_io_b2c_clk),
    .fpga_io_b2c_rst(clBridge_fpga_io_b2c_rst),
    .fpga_io_b2c_send(clBridge_fpga_io_b2c_send),
    .fpga_io_b2c_data(clBridge_fpga_io_b2c_data)
  );
  assign mem_axi4_0_awvalid = clBridge_io_master_awvalid; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_awid = clBridge_io_master_awid; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_awaddr = clBridge_io_master_awaddr; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_awlen = clBridge_io_master_awlen; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_awsize = clBridge_io_master_awsize; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_awburst = clBridge_io_master_awburst; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_wvalid = clBridge_io_master_wvalid; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_wdata = clBridge_io_master_wdata; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_wstrb = clBridge_io_master_wstrb; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_wlast = clBridge_io_master_wlast; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_bready = clBridge_io_master_bready; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_arvalid = clBridge_io_master_arvalid; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_arid = clBridge_io_master_arid; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_araddr = clBridge_io_master_araddr; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_arlen = clBridge_io_master_arlen; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_arsize = clBridge_io_master_arsize; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_arburst = clBridge_io_master_arburst; // @[TestHarness.scala 38:14]
  assign mem_axi4_0_rready = clBridge_io_master_rready; // @[TestHarness.scala 38:14]
  assign slave_axi4_mem_0_awready = clBridge_io_slave_awready; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_wready = clBridge_io_slave_wready; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_bvalid = clBridge_io_slave_bvalid; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_bid = clBridge_io_slave_bid; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_bresp = clBridge_io_slave_bresp; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_arready = clBridge_io_slave_arready; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_rvalid = clBridge_io_slave_rvalid; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_rid = clBridge_io_slave_rid; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_rdata = clBridge_io_slave_rdata; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_rresp = clBridge_io_slave_rresp; // @[TestHarness.scala 39:22]
  assign slave_axi4_mem_0_rlast = clBridge_io_slave_rlast; // @[TestHarness.scala 39:22]
  assign fpga_io_c2b_clk = clBridge_fpga_io_c2b_clk; // @[TestHarness.scala 40:11]
  assign fpga_io_c2b_rst = clBridge_fpga_io_c2b_rst; // @[TestHarness.scala 40:11]
  assign fpga_io_c2b_send = clBridge_fpga_io_c2b_send; // @[TestHarness.scala 40:11]
  assign fpga_io_c2b_data = clBridge_fpga_io_c2b_data; // @[TestHarness.scala 40:11]
  assign clBridge_clock = clock;
  assign clBridge_reset = reset;
  assign clBridge_io_master_awready = mem_axi4_0_awready; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_wready = mem_axi4_0_wready; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_bvalid = mem_axi4_0_bvalid; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_bid = mem_axi4_0_bid; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_bresp = mem_axi4_0_bresp; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_arready = mem_axi4_0_arready; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_rvalid = mem_axi4_0_rvalid; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_rid = mem_axi4_0_rid; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_rdata = mem_axi4_0_rdata; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_rresp = mem_axi4_0_rresp; // @[TestHarness.scala 38:14]
  assign clBridge_io_master_rlast = mem_axi4_0_rlast; // @[TestHarness.scala 38:14]
  assign clBridge_io_slave_awvalid = slave_axi4_mem_0_awvalid; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_awid = slave_axi4_mem_0_awid; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_awaddr = slave_axi4_mem_0_awaddr; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_awlen = slave_axi4_mem_0_awlen; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_awsize = slave_axi4_mem_0_awsize; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_awburst = slave_axi4_mem_0_awburst; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_wvalid = slave_axi4_mem_0_wvalid; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_wdata = slave_axi4_mem_0_wdata; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_wstrb = slave_axi4_mem_0_wstrb; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_wlast = slave_axi4_mem_0_wlast; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_bready = slave_axi4_mem_0_bready; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_arvalid = slave_axi4_mem_0_arvalid; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_arid = slave_axi4_mem_0_arid; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_araddr = slave_axi4_mem_0_araddr; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_arlen = slave_axi4_mem_0_arlen; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_arsize = slave_axi4_mem_0_arsize; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_arburst = slave_axi4_mem_0_arburst; // @[TestHarness.scala 39:22]
  assign clBridge_io_slave_rready = slave_axi4_mem_0_rready; // @[TestHarness.scala 39:22]
  assign clBridge_fpga_io_b2c_clk = fpga_io_b2c_clk; // @[TestHarness.scala 40:11]
  assign clBridge_fpga_io_b2c_rst = fpga_io_b2c_rst; // @[TestHarness.scala 40:11]
  assign clBridge_fpga_io_b2c_send = fpga_io_b2c_send; // @[TestHarness.scala 40:11]
  assign clBridge_fpga_io_b2c_data = fpga_io_b2c_data; // @[TestHarness.scala 40:11]
endmodule
module ram(
  input  [4:0]  R0_addr,
  input         R0_en,
  input         R0_clk,
  output [31:0] R0_data,
  input  [4:0]  W0_addr,
  input         W0_en,
  input         W0_clk,
  input  [31:0] W0_data
);
  wire [4:0] ram_ext_R0_addr;
  wire  ram_ext_R0_en;
  wire  ram_ext_R0_clk;
  wire [31:0] ram_ext_R0_data;
  wire [4:0] ram_ext_W0_addr;
  wire  ram_ext_W0_en;
  wire  ram_ext_W0_clk;
  wire [31:0] ram_ext_W0_data;
  ram_ext ram_ext (
    .R0_addr(ram_ext_R0_addr),
    .R0_en(ram_ext_R0_en),
    .R0_clk(ram_ext_R0_clk),
    .R0_data(ram_ext_R0_data),
    .W0_addr(ram_ext_W0_addr),
    .W0_en(ram_ext_W0_en),
    .W0_clk(ram_ext_W0_clk),
    .W0_data(ram_ext_W0_data)
  );
  assign ram_ext_R0_clk = R0_clk;
  assign ram_ext_R0_en = R0_en;
  assign ram_ext_R0_addr = R0_addr;
  assign R0_data = ram_ext_R0_data;
  assign ram_ext_W0_clk = W0_clk;
  assign ram_ext_W0_en = W0_en;
  assign ram_ext_W0_addr = W0_addr;
  assign ram_ext_W0_data = W0_data;
endmodule

module ram_ext(
  input W0_clk,
  input [4:0] W0_addr,
  input W0_en,
  input [31:0] W0_data,
  input R0_clk,
  input [4:0] R0_addr,
  input R0_en,
  output [31:0] R0_data
);

  reg reg_R0_ren;
  reg [4:0] reg_R0_addr;
  reg [31:0] ram [31:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 32; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
      reg_R0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge R0_clk)
    reg_R0_ren <= R0_en;
  always @(posedge R0_clk)
    if (R0_en) reg_R0_addr <= R0_addr;
  always @(posedge W0_clk)
    if (W0_en) begin
      ram[W0_addr][31:0] <= W0_data[31:0];
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] R0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      R0_random = {$random};
      reg_R0_ren = R0_random[0];
    end
  `endif
  always @(posedge R0_clk) R0_random <= {$random};
  assign R0_data = reg_R0_ren ? ram[reg_R0_addr] : R0_random[31:0];
  `else
  assign R0_data = ram[reg_R0_addr];
  `endif

endmodule
// See LICENSE.SiFive for license details.

//VCS coverage exclude_file

// No default parameter values are intended, nor does IEEE 1800-2012 require them (clause A.2.4 param_assignment),
// but Incisive demands them. These default values should never be used.
module plusarg_reader #(
   parameter FORMAT="borked=%d",
   parameter WIDTH=1,
   parameter [WIDTH-1:0] DEFAULT=0
) (
   output [WIDTH-1:0] out
);

`ifdef SYNTHESIS
assign out = DEFAULT;
`else
reg [WIDTH-1:0] myplus;
assign out = myplus;

initial begin
   if (!$value$plusargs(FORMAT, myplus)) myplus = DEFAULT;
end
`endif

endmodule
/* verilator lint_off UNOPTFLAT */

module EICG_wrapper(
  output out,
  input en,
  input test_en,
  input in
);

  reg en_latched /*verilator clock_enable*/;

  always @(*) begin
     if (!in) begin
        en_latched = en || test_en;
     end
  end

  assign out = en_latched && in;

endmodule
